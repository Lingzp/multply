$date
	Sat Jan 07 11:35:06 2023
$end
$version
	ModelSim Version 2020.1
$end
$timescale
	1ps
$end

$scope module Multiplier_Wrapper_tb $end
$var parameter 32 ! LIMIT $end
$var reg 1 " clock $end
$var reg 1 # reset $end
$var wire 1 $ m [63] $end
$var wire 1 % m [62] $end
$var wire 1 & m [61] $end
$var wire 1 ' m [60] $end
$var wire 1 ( m [59] $end
$var wire 1 ) m [58] $end
$var wire 1 * m [57] $end
$var wire 1 + m [56] $end
$var wire 1 , m [55] $end
$var wire 1 - m [54] $end
$var wire 1 . m [53] $end
$var wire 1 / m [52] $end
$var wire 1 0 m [51] $end
$var wire 1 1 m [50] $end
$var wire 1 2 m [49] $end
$var wire 1 3 m [48] $end
$var wire 1 4 m [47] $end
$var wire 1 5 m [46] $end
$var wire 1 6 m [45] $end
$var wire 1 7 m [44] $end
$var wire 1 8 m [43] $end
$var wire 1 9 m [42] $end
$var wire 1 : m [41] $end
$var wire 1 ; m [40] $end
$var wire 1 < m [39] $end
$var wire 1 = m [38] $end
$var wire 1 > m [37] $end
$var wire 1 ? m [36] $end
$var wire 1 @ m [35] $end
$var wire 1 A m [34] $end
$var wire 1 B m [33] $end
$var wire 1 C m [32] $end
$var wire 1 D m [31] $end
$var wire 1 E m [30] $end
$var wire 1 F m [29] $end
$var wire 1 G m [28] $end
$var wire 1 H m [27] $end
$var wire 1 I m [26] $end
$var wire 1 J m [25] $end
$var wire 1 K m [24] $end
$var wire 1 L m [23] $end
$var wire 1 M m [22] $end
$var wire 1 N m [21] $end
$var wire 1 O m [20] $end
$var wire 1 P m [19] $end
$var wire 1 Q m [18] $end
$var wire 1 R m [17] $end
$var wire 1 S m [16] $end
$var wire 1 T m [15] $end
$var wire 1 U m [14] $end
$var wire 1 V m [13] $end
$var wire 1 W m [12] $end
$var wire 1 X m [11] $end
$var wire 1 Y m [10] $end
$var wire 1 Z m [9] $end
$var wire 1 [ m [8] $end
$var wire 1 \ m [7] $end
$var wire 1 ] m [6] $end
$var wire 1 ^ m [5] $end
$var wire 1 _ m [4] $end
$var wire 1 ` m [3] $end
$var wire 1 a m [2] $end
$var wire 1 b m [1] $end
$var wire 1 c m [0] $end
$var reg 32 d a [31:0] $end
$var reg 32 e b [31:0] $end
$var wire 1 f golden_model [63] $end
$var wire 1 g golden_model [62] $end
$var wire 1 h golden_model [61] $end
$var wire 1 i golden_model [60] $end
$var wire 1 j golden_model [59] $end
$var wire 1 k golden_model [58] $end
$var wire 1 l golden_model [57] $end
$var wire 1 m golden_model [56] $end
$var wire 1 n golden_model [55] $end
$var wire 1 o golden_model [54] $end
$var wire 1 p golden_model [53] $end
$var wire 1 q golden_model [52] $end
$var wire 1 r golden_model [51] $end
$var wire 1 s golden_model [50] $end
$var wire 1 t golden_model [49] $end
$var wire 1 u golden_model [48] $end
$var wire 1 v golden_model [47] $end
$var wire 1 w golden_model [46] $end
$var wire 1 x golden_model [45] $end
$var wire 1 y golden_model [44] $end
$var wire 1 z golden_model [43] $end
$var wire 1 { golden_model [42] $end
$var wire 1 | golden_model [41] $end
$var wire 1 } golden_model [40] $end
$var wire 1 ~ golden_model [39] $end
$var wire 1 !! golden_model [38] $end
$var wire 1 "! golden_model [37] $end
$var wire 1 #! golden_model [36] $end
$var wire 1 $! golden_model [35] $end
$var wire 1 %! golden_model [34] $end
$var wire 1 &! golden_model [33] $end
$var wire 1 '! golden_model [32] $end
$var wire 1 (! golden_model [31] $end
$var wire 1 )! golden_model [30] $end
$var wire 1 *! golden_model [29] $end
$var wire 1 +! golden_model [28] $end
$var wire 1 ,! golden_model [27] $end
$var wire 1 -! golden_model [26] $end
$var wire 1 .! golden_model [25] $end
$var wire 1 /! golden_model [24] $end
$var wire 1 0! golden_model [23] $end
$var wire 1 1! golden_model [22] $end
$var wire 1 2! golden_model [21] $end
$var wire 1 3! golden_model [20] $end
$var wire 1 4! golden_model [19] $end
$var wire 1 5! golden_model [18] $end
$var wire 1 6! golden_model [17] $end
$var wire 1 7! golden_model [16] $end
$var wire 1 8! golden_model [15] $end
$var wire 1 9! golden_model [14] $end
$var wire 1 :! golden_model [13] $end
$var wire 1 ;! golden_model [12] $end
$var wire 1 <! golden_model [11] $end
$var wire 1 =! golden_model [10] $end
$var wire 1 >! golden_model [9] $end
$var wire 1 ?! golden_model [8] $end
$var wire 1 @! golden_model [7] $end
$var wire 1 A! golden_model [6] $end
$var wire 1 B! golden_model [5] $end
$var wire 1 C! golden_model [4] $end
$var wire 1 D! golden_model [3] $end
$var wire 1 E! golden_model [2] $end
$var wire 1 F! golden_model [1] $end
$var wire 1 G! golden_model [0] $end
$var reg 32 H! a_1p [31:0] $end
$var reg 32 I! b_1p [31:0] $end
$var reg 32 J! a_2p [31:0] $end
$var reg 32 K! b_2p [31:0] $end
$var reg 32 L! a_3p [31:0] $end
$var reg 32 M! b_3p [31:0] $end
$var reg 32 N! a_4p [31:0] $end
$var reg 32 O! b_4p [31:0] $end
$var reg 64 P! golden_model_1p [63:0] $end
$var reg 64 Q! golden_model_2p [63:0] $end
$var reg 64 R! golden_model_3p [63:0] $end
$var reg 64 S! golden_model_4p [63:0] $end

$scope module dut $end
$var wire 1 T! clk $end
$var wire 1 U! rst_n $end
$var wire 1 V! multiplicand [31] $end
$var wire 1 W! multiplicand [30] $end
$var wire 1 X! multiplicand [29] $end
$var wire 1 Y! multiplicand [28] $end
$var wire 1 Z! multiplicand [27] $end
$var wire 1 [! multiplicand [26] $end
$var wire 1 \! multiplicand [25] $end
$var wire 1 ]! multiplicand [24] $end
$var wire 1 ^! multiplicand [23] $end
$var wire 1 _! multiplicand [22] $end
$var wire 1 `! multiplicand [21] $end
$var wire 1 a! multiplicand [20] $end
$var wire 1 b! multiplicand [19] $end
$var wire 1 c! multiplicand [18] $end
$var wire 1 d! multiplicand [17] $end
$var wire 1 e! multiplicand [16] $end
$var wire 1 f! multiplicand [15] $end
$var wire 1 g! multiplicand [14] $end
$var wire 1 h! multiplicand [13] $end
$var wire 1 i! multiplicand [12] $end
$var wire 1 j! multiplicand [11] $end
$var wire 1 k! multiplicand [10] $end
$var wire 1 l! multiplicand [9] $end
$var wire 1 m! multiplicand [8] $end
$var wire 1 n! multiplicand [7] $end
$var wire 1 o! multiplicand [6] $end
$var wire 1 p! multiplicand [5] $end
$var wire 1 q! multiplicand [4] $end
$var wire 1 r! multiplicand [3] $end
$var wire 1 s! multiplicand [2] $end
$var wire 1 t! multiplicand [1] $end
$var wire 1 u! multiplicand [0] $end
$var wire 1 v! multiplier [31] $end
$var wire 1 w! multiplier [30] $end
$var wire 1 x! multiplier [29] $end
$var wire 1 y! multiplier [28] $end
$var wire 1 z! multiplier [27] $end
$var wire 1 {! multiplier [26] $end
$var wire 1 |! multiplier [25] $end
$var wire 1 }! multiplier [24] $end
$var wire 1 ~! multiplier [23] $end
$var wire 1 !" multiplier [22] $end
$var wire 1 "" multiplier [21] $end
$var wire 1 #" multiplier [20] $end
$var wire 1 $" multiplier [19] $end
$var wire 1 %" multiplier [18] $end
$var wire 1 &" multiplier [17] $end
$var wire 1 '" multiplier [16] $end
$var wire 1 (" multiplier [15] $end
$var wire 1 )" multiplier [14] $end
$var wire 1 *" multiplier [13] $end
$var wire 1 +" multiplier [12] $end
$var wire 1 ," multiplier [11] $end
$var wire 1 -" multiplier [10] $end
$var wire 1 ." multiplier [9] $end
$var wire 1 /" multiplier [8] $end
$var wire 1 0" multiplier [7] $end
$var wire 1 1" multiplier [6] $end
$var wire 1 2" multiplier [5] $end
$var wire 1 3" multiplier [4] $end
$var wire 1 4" multiplier [3] $end
$var wire 1 5" multiplier [2] $end
$var wire 1 6" multiplier [1] $end
$var wire 1 7" multiplier [0] $end
$var wire 1 $ product [63] $end
$var wire 1 % product [62] $end
$var wire 1 & product [61] $end
$var wire 1 ' product [60] $end
$var wire 1 ( product [59] $end
$var wire 1 ) product [58] $end
$var wire 1 * product [57] $end
$var wire 1 + product [56] $end
$var wire 1 , product [55] $end
$var wire 1 - product [54] $end
$var wire 1 . product [53] $end
$var wire 1 / product [52] $end
$var wire 1 0 product [51] $end
$var wire 1 1 product [50] $end
$var wire 1 2 product [49] $end
$var wire 1 3 product [48] $end
$var wire 1 4 product [47] $end
$var wire 1 5 product [46] $end
$var wire 1 6 product [45] $end
$var wire 1 7 product [44] $end
$var wire 1 8 product [43] $end
$var wire 1 9 product [42] $end
$var wire 1 : product [41] $end
$var wire 1 ; product [40] $end
$var wire 1 < product [39] $end
$var wire 1 = product [38] $end
$var wire 1 > product [37] $end
$var wire 1 ? product [36] $end
$var wire 1 @ product [35] $end
$var wire 1 A product [34] $end
$var wire 1 B product [33] $end
$var wire 1 C product [32] $end
$var wire 1 D product [31] $end
$var wire 1 E product [30] $end
$var wire 1 F product [29] $end
$var wire 1 G product [28] $end
$var wire 1 H product [27] $end
$var wire 1 I product [26] $end
$var wire 1 J product [25] $end
$var wire 1 K product [24] $end
$var wire 1 L product [23] $end
$var wire 1 M product [22] $end
$var wire 1 N product [21] $end
$var wire 1 O product [20] $end
$var wire 1 P product [19] $end
$var wire 1 Q product [18] $end
$var wire 1 R product [17] $end
$var wire 1 S product [16] $end
$var wire 1 T product [15] $end
$var wire 1 U product [14] $end
$var wire 1 V product [13] $end
$var wire 1 W product [12] $end
$var wire 1 X product [11] $end
$var wire 1 Y product [10] $end
$var wire 1 Z product [9] $end
$var wire 1 [ product [8] $end
$var wire 1 \ product [7] $end
$var wire 1 ] product [6] $end
$var wire 1 ^ product [5] $end
$var wire 1 _ product [4] $end
$var wire 1 ` product [3] $end
$var wire 1 a product [2] $end
$var wire 1 b product [1] $end
$var wire 1 c product [0] $end
$var wire 1 8" part_0 [32] $end
$var wire 1 9" part_0 [31] $end
$var wire 1 :" part_0 [30] $end
$var wire 1 ;" part_0 [29] $end
$var wire 1 <" part_0 [28] $end
$var wire 1 =" part_0 [27] $end
$var wire 1 >" part_0 [26] $end
$var wire 1 ?" part_0 [25] $end
$var wire 1 @" part_0 [24] $end
$var wire 1 A" part_0 [23] $end
$var wire 1 B" part_0 [22] $end
$var wire 1 C" part_0 [21] $end
$var wire 1 D" part_0 [20] $end
$var wire 1 E" part_0 [19] $end
$var wire 1 F" part_0 [18] $end
$var wire 1 G" part_0 [17] $end
$var wire 1 H" part_0 [16] $end
$var wire 1 I" part_0 [15] $end
$var wire 1 J" part_0 [14] $end
$var wire 1 K" part_0 [13] $end
$var wire 1 L" part_0 [12] $end
$var wire 1 M" part_0 [11] $end
$var wire 1 N" part_0 [10] $end
$var wire 1 O" part_0 [9] $end
$var wire 1 P" part_0 [8] $end
$var wire 1 Q" part_0 [7] $end
$var wire 1 R" part_0 [6] $end
$var wire 1 S" part_0 [5] $end
$var wire 1 T" part_0 [4] $end
$var wire 1 U" part_0 [3] $end
$var wire 1 V" part_0 [2] $end
$var wire 1 W" part_0 [1] $end
$var wire 1 X" part_0 [0] $end
$var wire 1 Y" part_1 [32] $end
$var wire 1 Z" part_1 [31] $end
$var wire 1 [" part_1 [30] $end
$var wire 1 \" part_1 [29] $end
$var wire 1 ]" part_1 [28] $end
$var wire 1 ^" part_1 [27] $end
$var wire 1 _" part_1 [26] $end
$var wire 1 `" part_1 [25] $end
$var wire 1 a" part_1 [24] $end
$var wire 1 b" part_1 [23] $end
$var wire 1 c" part_1 [22] $end
$var wire 1 d" part_1 [21] $end
$var wire 1 e" part_1 [20] $end
$var wire 1 f" part_1 [19] $end
$var wire 1 g" part_1 [18] $end
$var wire 1 h" part_1 [17] $end
$var wire 1 i" part_1 [16] $end
$var wire 1 j" part_1 [15] $end
$var wire 1 k" part_1 [14] $end
$var wire 1 l" part_1 [13] $end
$var wire 1 m" part_1 [12] $end
$var wire 1 n" part_1 [11] $end
$var wire 1 o" part_1 [10] $end
$var wire 1 p" part_1 [9] $end
$var wire 1 q" part_1 [8] $end
$var wire 1 r" part_1 [7] $end
$var wire 1 s" part_1 [6] $end
$var wire 1 t" part_1 [5] $end
$var wire 1 u" part_1 [4] $end
$var wire 1 v" part_1 [3] $end
$var wire 1 w" part_1 [2] $end
$var wire 1 x" part_1 [1] $end
$var wire 1 y" part_1 [0] $end
$var wire 1 z" part_2 [32] $end
$var wire 1 {" part_2 [31] $end
$var wire 1 |" part_2 [30] $end
$var wire 1 }" part_2 [29] $end
$var wire 1 ~" part_2 [28] $end
$var wire 1 !# part_2 [27] $end
$var wire 1 "# part_2 [26] $end
$var wire 1 ## part_2 [25] $end
$var wire 1 $# part_2 [24] $end
$var wire 1 %# part_2 [23] $end
$var wire 1 &# part_2 [22] $end
$var wire 1 '# part_2 [21] $end
$var wire 1 (# part_2 [20] $end
$var wire 1 )# part_2 [19] $end
$var wire 1 *# part_2 [18] $end
$var wire 1 +# part_2 [17] $end
$var wire 1 ,# part_2 [16] $end
$var wire 1 -# part_2 [15] $end
$var wire 1 .# part_2 [14] $end
$var wire 1 /# part_2 [13] $end
$var wire 1 0# part_2 [12] $end
$var wire 1 1# part_2 [11] $end
$var wire 1 2# part_2 [10] $end
$var wire 1 3# part_2 [9] $end
$var wire 1 4# part_2 [8] $end
$var wire 1 5# part_2 [7] $end
$var wire 1 6# part_2 [6] $end
$var wire 1 7# part_2 [5] $end
$var wire 1 8# part_2 [4] $end
$var wire 1 9# part_2 [3] $end
$var wire 1 :# part_2 [2] $end
$var wire 1 ;# part_2 [1] $end
$var wire 1 <# part_2 [0] $end
$var wire 1 =# part_3 [32] $end
$var wire 1 ># part_3 [31] $end
$var wire 1 ?# part_3 [30] $end
$var wire 1 @# part_3 [29] $end
$var wire 1 A# part_3 [28] $end
$var wire 1 B# part_3 [27] $end
$var wire 1 C# part_3 [26] $end
$var wire 1 D# part_3 [25] $end
$var wire 1 E# part_3 [24] $end
$var wire 1 F# part_3 [23] $end
$var wire 1 G# part_3 [22] $end
$var wire 1 H# part_3 [21] $end
$var wire 1 I# part_3 [20] $end
$var wire 1 J# part_3 [19] $end
$var wire 1 K# part_3 [18] $end
$var wire 1 L# part_3 [17] $end
$var wire 1 M# part_3 [16] $end
$var wire 1 N# part_3 [15] $end
$var wire 1 O# part_3 [14] $end
$var wire 1 P# part_3 [13] $end
$var wire 1 Q# part_3 [12] $end
$var wire 1 R# part_3 [11] $end
$var wire 1 S# part_3 [10] $end
$var wire 1 T# part_3 [9] $end
$var wire 1 U# part_3 [8] $end
$var wire 1 V# part_3 [7] $end
$var wire 1 W# part_3 [6] $end
$var wire 1 X# part_3 [5] $end
$var wire 1 Y# part_3 [4] $end
$var wire 1 Z# part_3 [3] $end
$var wire 1 [# part_3 [2] $end
$var wire 1 \# part_3 [1] $end
$var wire 1 ]# part_3 [0] $end
$var wire 1 ^# part_4 [32] $end
$var wire 1 _# part_4 [31] $end
$var wire 1 `# part_4 [30] $end
$var wire 1 a# part_4 [29] $end
$var wire 1 b# part_4 [28] $end
$var wire 1 c# part_4 [27] $end
$var wire 1 d# part_4 [26] $end
$var wire 1 e# part_4 [25] $end
$var wire 1 f# part_4 [24] $end
$var wire 1 g# part_4 [23] $end
$var wire 1 h# part_4 [22] $end
$var wire 1 i# part_4 [21] $end
$var wire 1 j# part_4 [20] $end
$var wire 1 k# part_4 [19] $end
$var wire 1 l# part_4 [18] $end
$var wire 1 m# part_4 [17] $end
$var wire 1 n# part_4 [16] $end
$var wire 1 o# part_4 [15] $end
$var wire 1 p# part_4 [14] $end
$var wire 1 q# part_4 [13] $end
$var wire 1 r# part_4 [12] $end
$var wire 1 s# part_4 [11] $end
$var wire 1 t# part_4 [10] $end
$var wire 1 u# part_4 [9] $end
$var wire 1 v# part_4 [8] $end
$var wire 1 w# part_4 [7] $end
$var wire 1 x# part_4 [6] $end
$var wire 1 y# part_4 [5] $end
$var wire 1 z# part_4 [4] $end
$var wire 1 {# part_4 [3] $end
$var wire 1 |# part_4 [2] $end
$var wire 1 }# part_4 [1] $end
$var wire 1 ~# part_4 [0] $end
$var wire 1 !$ part_5 [32] $end
$var wire 1 "$ part_5 [31] $end
$var wire 1 #$ part_5 [30] $end
$var wire 1 $$ part_5 [29] $end
$var wire 1 %$ part_5 [28] $end
$var wire 1 &$ part_5 [27] $end
$var wire 1 '$ part_5 [26] $end
$var wire 1 ($ part_5 [25] $end
$var wire 1 )$ part_5 [24] $end
$var wire 1 *$ part_5 [23] $end
$var wire 1 +$ part_5 [22] $end
$var wire 1 ,$ part_5 [21] $end
$var wire 1 -$ part_5 [20] $end
$var wire 1 .$ part_5 [19] $end
$var wire 1 /$ part_5 [18] $end
$var wire 1 0$ part_5 [17] $end
$var wire 1 1$ part_5 [16] $end
$var wire 1 2$ part_5 [15] $end
$var wire 1 3$ part_5 [14] $end
$var wire 1 4$ part_5 [13] $end
$var wire 1 5$ part_5 [12] $end
$var wire 1 6$ part_5 [11] $end
$var wire 1 7$ part_5 [10] $end
$var wire 1 8$ part_5 [9] $end
$var wire 1 9$ part_5 [8] $end
$var wire 1 :$ part_5 [7] $end
$var wire 1 ;$ part_5 [6] $end
$var wire 1 <$ part_5 [5] $end
$var wire 1 =$ part_5 [4] $end
$var wire 1 >$ part_5 [3] $end
$var wire 1 ?$ part_5 [2] $end
$var wire 1 @$ part_5 [1] $end
$var wire 1 A$ part_5 [0] $end
$var wire 1 B$ part_6 [32] $end
$var wire 1 C$ part_6 [31] $end
$var wire 1 D$ part_6 [30] $end
$var wire 1 E$ part_6 [29] $end
$var wire 1 F$ part_6 [28] $end
$var wire 1 G$ part_6 [27] $end
$var wire 1 H$ part_6 [26] $end
$var wire 1 I$ part_6 [25] $end
$var wire 1 J$ part_6 [24] $end
$var wire 1 K$ part_6 [23] $end
$var wire 1 L$ part_6 [22] $end
$var wire 1 M$ part_6 [21] $end
$var wire 1 N$ part_6 [20] $end
$var wire 1 O$ part_6 [19] $end
$var wire 1 P$ part_6 [18] $end
$var wire 1 Q$ part_6 [17] $end
$var wire 1 R$ part_6 [16] $end
$var wire 1 S$ part_6 [15] $end
$var wire 1 T$ part_6 [14] $end
$var wire 1 U$ part_6 [13] $end
$var wire 1 V$ part_6 [12] $end
$var wire 1 W$ part_6 [11] $end
$var wire 1 X$ part_6 [10] $end
$var wire 1 Y$ part_6 [9] $end
$var wire 1 Z$ part_6 [8] $end
$var wire 1 [$ part_6 [7] $end
$var wire 1 \$ part_6 [6] $end
$var wire 1 ]$ part_6 [5] $end
$var wire 1 ^$ part_6 [4] $end
$var wire 1 _$ part_6 [3] $end
$var wire 1 `$ part_6 [2] $end
$var wire 1 a$ part_6 [1] $end
$var wire 1 b$ part_6 [0] $end
$var wire 1 c$ part_7 [32] $end
$var wire 1 d$ part_7 [31] $end
$var wire 1 e$ part_7 [30] $end
$var wire 1 f$ part_7 [29] $end
$var wire 1 g$ part_7 [28] $end
$var wire 1 h$ part_7 [27] $end
$var wire 1 i$ part_7 [26] $end
$var wire 1 j$ part_7 [25] $end
$var wire 1 k$ part_7 [24] $end
$var wire 1 l$ part_7 [23] $end
$var wire 1 m$ part_7 [22] $end
$var wire 1 n$ part_7 [21] $end
$var wire 1 o$ part_7 [20] $end
$var wire 1 p$ part_7 [19] $end
$var wire 1 q$ part_7 [18] $end
$var wire 1 r$ part_7 [17] $end
$var wire 1 s$ part_7 [16] $end
$var wire 1 t$ part_7 [15] $end
$var wire 1 u$ part_7 [14] $end
$var wire 1 v$ part_7 [13] $end
$var wire 1 w$ part_7 [12] $end
$var wire 1 x$ part_7 [11] $end
$var wire 1 y$ part_7 [10] $end
$var wire 1 z$ part_7 [9] $end
$var wire 1 {$ part_7 [8] $end
$var wire 1 |$ part_7 [7] $end
$var wire 1 }$ part_7 [6] $end
$var wire 1 ~$ part_7 [5] $end
$var wire 1 !% part_7 [4] $end
$var wire 1 "% part_7 [3] $end
$var wire 1 #% part_7 [2] $end
$var wire 1 $% part_7 [1] $end
$var wire 1 %% part_7 [0] $end
$var wire 1 &% part_8 [32] $end
$var wire 1 '% part_8 [31] $end
$var wire 1 (% part_8 [30] $end
$var wire 1 )% part_8 [29] $end
$var wire 1 *% part_8 [28] $end
$var wire 1 +% part_8 [27] $end
$var wire 1 ,% part_8 [26] $end
$var wire 1 -% part_8 [25] $end
$var wire 1 .% part_8 [24] $end
$var wire 1 /% part_8 [23] $end
$var wire 1 0% part_8 [22] $end
$var wire 1 1% part_8 [21] $end
$var wire 1 2% part_8 [20] $end
$var wire 1 3% part_8 [19] $end
$var wire 1 4% part_8 [18] $end
$var wire 1 5% part_8 [17] $end
$var wire 1 6% part_8 [16] $end
$var wire 1 7% part_8 [15] $end
$var wire 1 8% part_8 [14] $end
$var wire 1 9% part_8 [13] $end
$var wire 1 :% part_8 [12] $end
$var wire 1 ;% part_8 [11] $end
$var wire 1 <% part_8 [10] $end
$var wire 1 =% part_8 [9] $end
$var wire 1 >% part_8 [8] $end
$var wire 1 ?% part_8 [7] $end
$var wire 1 @% part_8 [6] $end
$var wire 1 A% part_8 [5] $end
$var wire 1 B% part_8 [4] $end
$var wire 1 C% part_8 [3] $end
$var wire 1 D% part_8 [2] $end
$var wire 1 E% part_8 [1] $end
$var wire 1 F% part_8 [0] $end
$var wire 1 G% part_9 [32] $end
$var wire 1 H% part_9 [31] $end
$var wire 1 I% part_9 [30] $end
$var wire 1 J% part_9 [29] $end
$var wire 1 K% part_9 [28] $end
$var wire 1 L% part_9 [27] $end
$var wire 1 M% part_9 [26] $end
$var wire 1 N% part_9 [25] $end
$var wire 1 O% part_9 [24] $end
$var wire 1 P% part_9 [23] $end
$var wire 1 Q% part_9 [22] $end
$var wire 1 R% part_9 [21] $end
$var wire 1 S% part_9 [20] $end
$var wire 1 T% part_9 [19] $end
$var wire 1 U% part_9 [18] $end
$var wire 1 V% part_9 [17] $end
$var wire 1 W% part_9 [16] $end
$var wire 1 X% part_9 [15] $end
$var wire 1 Y% part_9 [14] $end
$var wire 1 Z% part_9 [13] $end
$var wire 1 [% part_9 [12] $end
$var wire 1 \% part_9 [11] $end
$var wire 1 ]% part_9 [10] $end
$var wire 1 ^% part_9 [9] $end
$var wire 1 _% part_9 [8] $end
$var wire 1 `% part_9 [7] $end
$var wire 1 a% part_9 [6] $end
$var wire 1 b% part_9 [5] $end
$var wire 1 c% part_9 [4] $end
$var wire 1 d% part_9 [3] $end
$var wire 1 e% part_9 [2] $end
$var wire 1 f% part_9 [1] $end
$var wire 1 g% part_9 [0] $end
$var wire 1 h% part_10 [32] $end
$var wire 1 i% part_10 [31] $end
$var wire 1 j% part_10 [30] $end
$var wire 1 k% part_10 [29] $end
$var wire 1 l% part_10 [28] $end
$var wire 1 m% part_10 [27] $end
$var wire 1 n% part_10 [26] $end
$var wire 1 o% part_10 [25] $end
$var wire 1 p% part_10 [24] $end
$var wire 1 q% part_10 [23] $end
$var wire 1 r% part_10 [22] $end
$var wire 1 s% part_10 [21] $end
$var wire 1 t% part_10 [20] $end
$var wire 1 u% part_10 [19] $end
$var wire 1 v% part_10 [18] $end
$var wire 1 w% part_10 [17] $end
$var wire 1 x% part_10 [16] $end
$var wire 1 y% part_10 [15] $end
$var wire 1 z% part_10 [14] $end
$var wire 1 {% part_10 [13] $end
$var wire 1 |% part_10 [12] $end
$var wire 1 }% part_10 [11] $end
$var wire 1 ~% part_10 [10] $end
$var wire 1 !& part_10 [9] $end
$var wire 1 "& part_10 [8] $end
$var wire 1 #& part_10 [7] $end
$var wire 1 $& part_10 [6] $end
$var wire 1 %& part_10 [5] $end
$var wire 1 && part_10 [4] $end
$var wire 1 '& part_10 [3] $end
$var wire 1 (& part_10 [2] $end
$var wire 1 )& part_10 [1] $end
$var wire 1 *& part_10 [0] $end
$var wire 1 +& part_11 [32] $end
$var wire 1 ,& part_11 [31] $end
$var wire 1 -& part_11 [30] $end
$var wire 1 .& part_11 [29] $end
$var wire 1 /& part_11 [28] $end
$var wire 1 0& part_11 [27] $end
$var wire 1 1& part_11 [26] $end
$var wire 1 2& part_11 [25] $end
$var wire 1 3& part_11 [24] $end
$var wire 1 4& part_11 [23] $end
$var wire 1 5& part_11 [22] $end
$var wire 1 6& part_11 [21] $end
$var wire 1 7& part_11 [20] $end
$var wire 1 8& part_11 [19] $end
$var wire 1 9& part_11 [18] $end
$var wire 1 :& part_11 [17] $end
$var wire 1 ;& part_11 [16] $end
$var wire 1 <& part_11 [15] $end
$var wire 1 =& part_11 [14] $end
$var wire 1 >& part_11 [13] $end
$var wire 1 ?& part_11 [12] $end
$var wire 1 @& part_11 [11] $end
$var wire 1 A& part_11 [10] $end
$var wire 1 B& part_11 [9] $end
$var wire 1 C& part_11 [8] $end
$var wire 1 D& part_11 [7] $end
$var wire 1 E& part_11 [6] $end
$var wire 1 F& part_11 [5] $end
$var wire 1 G& part_11 [4] $end
$var wire 1 H& part_11 [3] $end
$var wire 1 I& part_11 [2] $end
$var wire 1 J& part_11 [1] $end
$var wire 1 K& part_11 [0] $end
$var wire 1 L& part_12 [32] $end
$var wire 1 M& part_12 [31] $end
$var wire 1 N& part_12 [30] $end
$var wire 1 O& part_12 [29] $end
$var wire 1 P& part_12 [28] $end
$var wire 1 Q& part_12 [27] $end
$var wire 1 R& part_12 [26] $end
$var wire 1 S& part_12 [25] $end
$var wire 1 T& part_12 [24] $end
$var wire 1 U& part_12 [23] $end
$var wire 1 V& part_12 [22] $end
$var wire 1 W& part_12 [21] $end
$var wire 1 X& part_12 [20] $end
$var wire 1 Y& part_12 [19] $end
$var wire 1 Z& part_12 [18] $end
$var wire 1 [& part_12 [17] $end
$var wire 1 \& part_12 [16] $end
$var wire 1 ]& part_12 [15] $end
$var wire 1 ^& part_12 [14] $end
$var wire 1 _& part_12 [13] $end
$var wire 1 `& part_12 [12] $end
$var wire 1 a& part_12 [11] $end
$var wire 1 b& part_12 [10] $end
$var wire 1 c& part_12 [9] $end
$var wire 1 d& part_12 [8] $end
$var wire 1 e& part_12 [7] $end
$var wire 1 f& part_12 [6] $end
$var wire 1 g& part_12 [5] $end
$var wire 1 h& part_12 [4] $end
$var wire 1 i& part_12 [3] $end
$var wire 1 j& part_12 [2] $end
$var wire 1 k& part_12 [1] $end
$var wire 1 l& part_12 [0] $end
$var wire 1 m& part_13 [32] $end
$var wire 1 n& part_13 [31] $end
$var wire 1 o& part_13 [30] $end
$var wire 1 p& part_13 [29] $end
$var wire 1 q& part_13 [28] $end
$var wire 1 r& part_13 [27] $end
$var wire 1 s& part_13 [26] $end
$var wire 1 t& part_13 [25] $end
$var wire 1 u& part_13 [24] $end
$var wire 1 v& part_13 [23] $end
$var wire 1 w& part_13 [22] $end
$var wire 1 x& part_13 [21] $end
$var wire 1 y& part_13 [20] $end
$var wire 1 z& part_13 [19] $end
$var wire 1 {& part_13 [18] $end
$var wire 1 |& part_13 [17] $end
$var wire 1 }& part_13 [16] $end
$var wire 1 ~& part_13 [15] $end
$var wire 1 !' part_13 [14] $end
$var wire 1 "' part_13 [13] $end
$var wire 1 #' part_13 [12] $end
$var wire 1 $' part_13 [11] $end
$var wire 1 %' part_13 [10] $end
$var wire 1 &' part_13 [9] $end
$var wire 1 '' part_13 [8] $end
$var wire 1 (' part_13 [7] $end
$var wire 1 )' part_13 [6] $end
$var wire 1 *' part_13 [5] $end
$var wire 1 +' part_13 [4] $end
$var wire 1 ,' part_13 [3] $end
$var wire 1 -' part_13 [2] $end
$var wire 1 .' part_13 [1] $end
$var wire 1 /' part_13 [0] $end
$var wire 1 0' part_14 [32] $end
$var wire 1 1' part_14 [31] $end
$var wire 1 2' part_14 [30] $end
$var wire 1 3' part_14 [29] $end
$var wire 1 4' part_14 [28] $end
$var wire 1 5' part_14 [27] $end
$var wire 1 6' part_14 [26] $end
$var wire 1 7' part_14 [25] $end
$var wire 1 8' part_14 [24] $end
$var wire 1 9' part_14 [23] $end
$var wire 1 :' part_14 [22] $end
$var wire 1 ;' part_14 [21] $end
$var wire 1 <' part_14 [20] $end
$var wire 1 =' part_14 [19] $end
$var wire 1 >' part_14 [18] $end
$var wire 1 ?' part_14 [17] $end
$var wire 1 @' part_14 [16] $end
$var wire 1 A' part_14 [15] $end
$var wire 1 B' part_14 [14] $end
$var wire 1 C' part_14 [13] $end
$var wire 1 D' part_14 [12] $end
$var wire 1 E' part_14 [11] $end
$var wire 1 F' part_14 [10] $end
$var wire 1 G' part_14 [9] $end
$var wire 1 H' part_14 [8] $end
$var wire 1 I' part_14 [7] $end
$var wire 1 J' part_14 [6] $end
$var wire 1 K' part_14 [5] $end
$var wire 1 L' part_14 [4] $end
$var wire 1 M' part_14 [3] $end
$var wire 1 N' part_14 [2] $end
$var wire 1 O' part_14 [1] $end
$var wire 1 P' part_14 [0] $end
$var wire 1 Q' part_15 [32] $end
$var wire 1 R' part_15 [31] $end
$var wire 1 S' part_15 [30] $end
$var wire 1 T' part_15 [29] $end
$var wire 1 U' part_15 [28] $end
$var wire 1 V' part_15 [27] $end
$var wire 1 W' part_15 [26] $end
$var wire 1 X' part_15 [25] $end
$var wire 1 Y' part_15 [24] $end
$var wire 1 Z' part_15 [23] $end
$var wire 1 [' part_15 [22] $end
$var wire 1 \' part_15 [21] $end
$var wire 1 ]' part_15 [20] $end
$var wire 1 ^' part_15 [19] $end
$var wire 1 _' part_15 [18] $end
$var wire 1 `' part_15 [17] $end
$var wire 1 a' part_15 [16] $end
$var wire 1 b' part_15 [15] $end
$var wire 1 c' part_15 [14] $end
$var wire 1 d' part_15 [13] $end
$var wire 1 e' part_15 [12] $end
$var wire 1 f' part_15 [11] $end
$var wire 1 g' part_15 [10] $end
$var wire 1 h' part_15 [9] $end
$var wire 1 i' part_15 [8] $end
$var wire 1 j' part_15 [7] $end
$var wire 1 k' part_15 [6] $end
$var wire 1 l' part_15 [5] $end
$var wire 1 m' part_15 [4] $end
$var wire 1 n' part_15 [3] $end
$var wire 1 o' part_15 [2] $end
$var wire 1 p' part_15 [1] $end
$var wire 1 q' part_15 [0] $end
$var wire 1 r' part_16 [30] $end
$var wire 1 s' part_16 [29] $end
$var wire 1 t' part_16 [28] $end
$var wire 1 u' part_16 [27] $end
$var wire 1 v' part_16 [26] $end
$var wire 1 w' part_16 [25] $end
$var wire 1 x' part_16 [24] $end
$var wire 1 y' part_16 [23] $end
$var wire 1 z' part_16 [22] $end
$var wire 1 {' part_16 [21] $end
$var wire 1 |' part_16 [20] $end
$var wire 1 }' part_16 [19] $end
$var wire 1 ~' part_16 [18] $end
$var wire 1 !( part_16 [17] $end
$var wire 1 "( part_16 [16] $end
$var wire 1 #( part_16 [15] $end
$var wire 1 $( part_16 [14] $end
$var wire 1 %( part_16 [13] $end
$var wire 1 &( part_16 [12] $end
$var wire 1 '( part_16 [11] $end
$var wire 1 (( part_16 [10] $end
$var wire 1 )( part_16 [9] $end
$var wire 1 *( part_16 [8] $end
$var wire 1 +( part_16 [7] $end
$var wire 1 ,( part_16 [6] $end
$var wire 1 -( part_16 [5] $end
$var wire 1 .( part_16 [4] $end
$var wire 1 /( part_16 [3] $end
$var wire 1 0( part_16 [2] $end
$var wire 1 1( part_16 [1] $end
$var wire 1 2( part_16 [0] $end
$var wire 1 3( h0 [1] $end
$var wire 1 4( h0 [0] $end
$var wire 1 5( h1 [1] $end
$var wire 1 6( h1 [0] $end
$var wire 1 7( h2 [1] $end
$var wire 1 8( h2 [0] $end
$var wire 1 9( h3 [1] $end
$var wire 1 :( h3 [0] $end
$var wire 1 ;( h4 [1] $end
$var wire 1 <( h4 [0] $end
$var wire 1 =( h5 [1] $end
$var wire 1 >( h5 [0] $end
$var wire 1 ?( h6 [1] $end
$var wire 1 @( h6 [0] $end
$var wire 1 A( h7 [1] $end
$var wire 1 B( h7 [0] $end
$var wire 1 C( h8 [1] $end
$var wire 1 D( h8 [0] $end
$var wire 1 E( h9 [1] $end
$var wire 1 F( h9 [0] $end
$var wire 1 G( h10 [1] $end
$var wire 1 H( h10 [0] $end
$var wire 1 I( h11 [1] $end
$var wire 1 J( h11 [0] $end
$var wire 1 K( h12 [1] $end
$var wire 1 L( h12 [0] $end
$var wire 1 M( h13 [1] $end
$var wire 1 N( h13 [0] $end
$var wire 1 O( h14 [1] $end
$var wire 1 P( h14 [0] $end
$var wire 1 Q( h15 [1] $end
$var wire 1 R( h15 [0] $end
$var wire 1 S( multiplicand_not [31] $end
$var wire 1 T( multiplicand_not [30] $end
$var wire 1 U( multiplicand_not [29] $end
$var wire 1 V( multiplicand_not [28] $end
$var wire 1 W( multiplicand_not [27] $end
$var wire 1 X( multiplicand_not [26] $end
$var wire 1 Y( multiplicand_not [25] $end
$var wire 1 Z( multiplicand_not [24] $end
$var wire 1 [( multiplicand_not [23] $end
$var wire 1 \( multiplicand_not [22] $end
$var wire 1 ]( multiplicand_not [21] $end
$var wire 1 ^( multiplicand_not [20] $end
$var wire 1 _( multiplicand_not [19] $end
$var wire 1 `( multiplicand_not [18] $end
$var wire 1 a( multiplicand_not [17] $end
$var wire 1 b( multiplicand_not [16] $end
$var wire 1 c( multiplicand_not [15] $end
$var wire 1 d( multiplicand_not [14] $end
$var wire 1 e( multiplicand_not [13] $end
$var wire 1 f( multiplicand_not [12] $end
$var wire 1 g( multiplicand_not [11] $end
$var wire 1 h( multiplicand_not [10] $end
$var wire 1 i( multiplicand_not [9] $end
$var wire 1 j( multiplicand_not [8] $end
$var wire 1 k( multiplicand_not [7] $end
$var wire 1 l( multiplicand_not [6] $end
$var wire 1 m( multiplicand_not [5] $end
$var wire 1 n( multiplicand_not [4] $end
$var wire 1 o( multiplicand_not [3] $end
$var wire 1 p( multiplicand_not [2] $end
$var wire 1 q( multiplicand_not [1] $end
$var wire 1 r( multiplicand_not [0] $end
$var wire 1 s( sign [16] $end
$var wire 1 t( sign [15] $end
$var wire 1 u( sign [14] $end
$var wire 1 v( sign [13] $end
$var wire 1 w( sign [12] $end
$var wire 1 x( sign [11] $end
$var wire 1 y( sign [10] $end
$var wire 1 z( sign [9] $end
$var wire 1 {( sign [8] $end
$var wire 1 |( sign [7] $end
$var wire 1 }( sign [6] $end
$var wire 1 ~( sign [5] $end
$var wire 1 !) sign [4] $end
$var wire 1 ") sign [3] $end
$var wire 1 #) sign [2] $end
$var wire 1 $) sign [1] $end
$var wire 1 %) sign [0] $end
$var wire 1 &) l1_1_0 [35] $end
$var wire 1 ') l1_1_0 [34] $end
$var wire 1 () l1_1_0 [33] $end
$var wire 1 )) l1_1_0 [32] $end
$var wire 1 *) l1_1_0 [31] $end
$var wire 1 +) l1_1_0 [30] $end
$var wire 1 ,) l1_1_0 [29] $end
$var wire 1 -) l1_1_0 [28] $end
$var wire 1 .) l1_1_0 [27] $end
$var wire 1 /) l1_1_0 [26] $end
$var wire 1 0) l1_1_0 [25] $end
$var wire 1 1) l1_1_0 [24] $end
$var wire 1 2) l1_1_0 [23] $end
$var wire 1 3) l1_1_0 [22] $end
$var wire 1 4) l1_1_0 [21] $end
$var wire 1 5) l1_1_0 [20] $end
$var wire 1 6) l1_1_0 [19] $end
$var wire 1 7) l1_1_0 [18] $end
$var wire 1 8) l1_1_0 [17] $end
$var wire 1 9) l1_1_0 [16] $end
$var wire 1 :) l1_1_0 [15] $end
$var wire 1 ;) l1_1_0 [14] $end
$var wire 1 <) l1_1_0 [13] $end
$var wire 1 =) l1_1_0 [12] $end
$var wire 1 >) l1_1_0 [11] $end
$var wire 1 ?) l1_1_0 [10] $end
$var wire 1 @) l1_1_0 [9] $end
$var wire 1 A) l1_1_0 [8] $end
$var wire 1 B) l1_1_0 [7] $end
$var wire 1 C) l1_1_0 [6] $end
$var wire 1 D) l1_1_0 [5] $end
$var wire 1 E) l1_1_0 [4] $end
$var wire 1 F) l1_1_0 [3] $end
$var wire 1 G) l1_1_0 [2] $end
$var wire 1 H) l1_1_0 [1] $end
$var wire 1 I) l1_1_0 [0] $end
$var wire 1 J) l1_1_1 [35] $end
$var wire 1 K) l1_1_1 [34] $end
$var wire 1 L) l1_1_1 [33] $end
$var wire 1 M) l1_1_1 [32] $end
$var wire 1 N) l1_1_1 [31] $end
$var wire 1 O) l1_1_1 [30] $end
$var wire 1 P) l1_1_1 [29] $end
$var wire 1 Q) l1_1_1 [28] $end
$var wire 1 R) l1_1_1 [27] $end
$var wire 1 S) l1_1_1 [26] $end
$var wire 1 T) l1_1_1 [25] $end
$var wire 1 U) l1_1_1 [24] $end
$var wire 1 V) l1_1_1 [23] $end
$var wire 1 W) l1_1_1 [22] $end
$var wire 1 X) l1_1_1 [21] $end
$var wire 1 Y) l1_1_1 [20] $end
$var wire 1 Z) l1_1_1 [19] $end
$var wire 1 [) l1_1_1 [18] $end
$var wire 1 \) l1_1_1 [17] $end
$var wire 1 ]) l1_1_1 [16] $end
$var wire 1 ^) l1_1_1 [15] $end
$var wire 1 _) l1_1_1 [14] $end
$var wire 1 `) l1_1_1 [13] $end
$var wire 1 a) l1_1_1 [12] $end
$var wire 1 b) l1_1_1 [11] $end
$var wire 1 c) l1_1_1 [10] $end
$var wire 1 d) l1_1_1 [9] $end
$var wire 1 e) l1_1_1 [8] $end
$var wire 1 f) l1_1_1 [7] $end
$var wire 1 g) l1_1_1 [6] $end
$var wire 1 h) l1_1_1 [5] $end
$var wire 1 i) l1_1_1 [4] $end
$var wire 1 j) l1_1_1 [3] $end
$var wire 1 k) l1_1_1 [2] $end
$var wire 1 l) l1_1_1 [1] $end
$var wire 1 m) l1_1_1 [0] $end
$var wire 1 n) l1_1_2 [35] $end
$var wire 1 o) l1_1_2 [34] $end
$var wire 1 p) l1_1_2 [33] $end
$var wire 1 q) l1_1_2 [32] $end
$var wire 1 r) l1_1_2 [31] $end
$var wire 1 s) l1_1_2 [30] $end
$var wire 1 t) l1_1_2 [29] $end
$var wire 1 u) l1_1_2 [28] $end
$var wire 1 v) l1_1_2 [27] $end
$var wire 1 w) l1_1_2 [26] $end
$var wire 1 x) l1_1_2 [25] $end
$var wire 1 y) l1_1_2 [24] $end
$var wire 1 z) l1_1_2 [23] $end
$var wire 1 {) l1_1_2 [22] $end
$var wire 1 |) l1_1_2 [21] $end
$var wire 1 }) l1_1_2 [20] $end
$var wire 1 ~) l1_1_2 [19] $end
$var wire 1 !* l1_1_2 [18] $end
$var wire 1 "* l1_1_2 [17] $end
$var wire 1 #* l1_1_2 [16] $end
$var wire 1 $* l1_1_2 [15] $end
$var wire 1 %* l1_1_2 [14] $end
$var wire 1 &* l1_1_2 [13] $end
$var wire 1 '* l1_1_2 [12] $end
$var wire 1 (* l1_1_2 [11] $end
$var wire 1 )* l1_1_2 [10] $end
$var wire 1 ** l1_1_2 [9] $end
$var wire 1 +* l1_1_2 [8] $end
$var wire 1 ,* l1_1_2 [7] $end
$var wire 1 -* l1_1_2 [6] $end
$var wire 1 .* l1_1_2 [5] $end
$var wire 1 /* l1_1_2 [4] $end
$var wire 1 0* l1_1_2 [3] $end
$var wire 1 1* l1_1_2 [2] $end
$var wire 1 2* l1_1_2 [1] $end
$var wire 1 3* l1_1_2 [0] $end
$var wire 1 4* l1_1_cin [35] $end
$var wire 1 5* l1_1_cin [34] $end
$var wire 1 6* l1_1_cin [33] $end
$var wire 1 7* l1_1_cin [32] $end
$var wire 1 8* l1_1_cin [31] $end
$var wire 1 9* l1_1_cin [30] $end
$var wire 1 :* l1_1_cin [29] $end
$var wire 1 ;* l1_1_cin [28] $end
$var wire 1 <* l1_1_cin [27] $end
$var wire 1 =* l1_1_cin [26] $end
$var wire 1 >* l1_1_cin [25] $end
$var wire 1 ?* l1_1_cin [24] $end
$var wire 1 @* l1_1_cin [23] $end
$var wire 1 A* l1_1_cin [22] $end
$var wire 1 B* l1_1_cin [21] $end
$var wire 1 C* l1_1_cin [20] $end
$var wire 1 D* l1_1_cin [19] $end
$var wire 1 E* l1_1_cin [18] $end
$var wire 1 F* l1_1_cin [17] $end
$var wire 1 G* l1_1_cin [16] $end
$var wire 1 H* l1_1_cin [15] $end
$var wire 1 I* l1_1_cin [14] $end
$var wire 1 J* l1_1_cin [13] $end
$var wire 1 K* l1_1_cin [12] $end
$var wire 1 L* l1_1_cin [11] $end
$var wire 1 M* l1_1_cin [10] $end
$var wire 1 N* l1_1_cin [9] $end
$var wire 1 O* l1_1_cin [8] $end
$var wire 1 P* l1_1_cin [7] $end
$var wire 1 Q* l1_1_cin [6] $end
$var wire 1 R* l1_1_cin [5] $end
$var wire 1 S* l1_1_cin [4] $end
$var wire 1 T* l1_1_cin [3] $end
$var wire 1 U* l1_1_cin [2] $end
$var wire 1 V* l1_1_cin [1] $end
$var wire 1 W* l1_1_cin [0] $end
$var wire 1 X* l1_1_cout [35] $end
$var wire 1 Y* l1_1_cout [34] $end
$var wire 1 Z* l1_1_cout [33] $end
$var wire 1 [* l1_1_cout [32] $end
$var wire 1 \* l1_1_cout [31] $end
$var wire 1 ]* l1_1_cout [30] $end
$var wire 1 ^* l1_1_cout [29] $end
$var wire 1 _* l1_1_cout [28] $end
$var wire 1 `* l1_1_cout [27] $end
$var wire 1 a* l1_1_cout [26] $end
$var wire 1 b* l1_1_cout [25] $end
$var wire 1 c* l1_1_cout [24] $end
$var wire 1 d* l1_1_cout [23] $end
$var wire 1 e* l1_1_cout [22] $end
$var wire 1 f* l1_1_cout [21] $end
$var wire 1 g* l1_1_cout [20] $end
$var wire 1 h* l1_1_cout [19] $end
$var wire 1 i* l1_1_cout [18] $end
$var wire 1 j* l1_1_cout [17] $end
$var wire 1 k* l1_1_cout [16] $end
$var wire 1 l* l1_1_cout [15] $end
$var wire 1 m* l1_1_cout [14] $end
$var wire 1 n* l1_1_cout [13] $end
$var wire 1 o* l1_1_cout [12] $end
$var wire 1 p* l1_1_cout [11] $end
$var wire 1 q* l1_1_cout [10] $end
$var wire 1 r* l1_1_cout [9] $end
$var wire 1 s* l1_1_cout [8] $end
$var wire 1 t* l1_1_cout [7] $end
$var wire 1 u* l1_1_cout [6] $end
$var wire 1 v* l1_1_cout [5] $end
$var wire 1 w* l1_1_cout [4] $end
$var wire 1 x* l1_1_cout [3] $end
$var wire 1 y* l1_1_cout [2] $end
$var wire 1 z* l1_1_cout [1] $end
$var wire 1 {* l1_1_cout [0] $end
$var wire 1 |* l1_1_s [35] $end
$var wire 1 }* l1_1_s [34] $end
$var wire 1 ~* l1_1_s [33] $end
$var wire 1 !+ l1_1_s [32] $end
$var wire 1 "+ l1_1_s [31] $end
$var wire 1 #+ l1_1_s [30] $end
$var wire 1 $+ l1_1_s [29] $end
$var wire 1 %+ l1_1_s [28] $end
$var wire 1 &+ l1_1_s [27] $end
$var wire 1 '+ l1_1_s [26] $end
$var wire 1 (+ l1_1_s [25] $end
$var wire 1 )+ l1_1_s [24] $end
$var wire 1 *+ l1_1_s [23] $end
$var wire 1 ++ l1_1_s [22] $end
$var wire 1 ,+ l1_1_s [21] $end
$var wire 1 -+ l1_1_s [20] $end
$var wire 1 .+ l1_1_s [19] $end
$var wire 1 /+ l1_1_s [18] $end
$var wire 1 0+ l1_1_s [17] $end
$var wire 1 1+ l1_1_s [16] $end
$var wire 1 2+ l1_1_s [15] $end
$var wire 1 3+ l1_1_s [14] $end
$var wire 1 4+ l1_1_s [13] $end
$var wire 1 5+ l1_1_s [12] $end
$var wire 1 6+ l1_1_s [11] $end
$var wire 1 7+ l1_1_s [10] $end
$var wire 1 8+ l1_1_s [9] $end
$var wire 1 9+ l1_1_s [8] $end
$var wire 1 :+ l1_1_s [7] $end
$var wire 1 ;+ l1_1_s [6] $end
$var wire 1 <+ l1_1_s [5] $end
$var wire 1 =+ l1_1_s [4] $end
$var wire 1 >+ l1_1_s [3] $end
$var wire 1 ?+ l1_1_s [2] $end
$var wire 1 @+ l1_1_s [1] $end
$var wire 1 A+ l1_1_s [0] $end
$var wire 1 B+ l1_1_ca [35] $end
$var wire 1 C+ l1_1_ca [34] $end
$var wire 1 D+ l1_1_ca [33] $end
$var wire 1 E+ l1_1_ca [32] $end
$var wire 1 F+ l1_1_ca [31] $end
$var wire 1 G+ l1_1_ca [30] $end
$var wire 1 H+ l1_1_ca [29] $end
$var wire 1 I+ l1_1_ca [28] $end
$var wire 1 J+ l1_1_ca [27] $end
$var wire 1 K+ l1_1_ca [26] $end
$var wire 1 L+ l1_1_ca [25] $end
$var wire 1 M+ l1_1_ca [24] $end
$var wire 1 N+ l1_1_ca [23] $end
$var wire 1 O+ l1_1_ca [22] $end
$var wire 1 P+ l1_1_ca [21] $end
$var wire 1 Q+ l1_1_ca [20] $end
$var wire 1 R+ l1_1_ca [19] $end
$var wire 1 S+ l1_1_ca [18] $end
$var wire 1 T+ l1_1_ca [17] $end
$var wire 1 U+ l1_1_ca [16] $end
$var wire 1 V+ l1_1_ca [15] $end
$var wire 1 W+ l1_1_ca [14] $end
$var wire 1 X+ l1_1_ca [13] $end
$var wire 1 Y+ l1_1_ca [12] $end
$var wire 1 Z+ l1_1_ca [11] $end
$var wire 1 [+ l1_1_ca [10] $end
$var wire 1 \+ l1_1_ca [9] $end
$var wire 1 ]+ l1_1_ca [8] $end
$var wire 1 ^+ l1_1_ca [7] $end
$var wire 1 _+ l1_1_ca [6] $end
$var wire 1 `+ l1_1_ca [5] $end
$var wire 1 a+ l1_1_ca [4] $end
$var wire 1 b+ l1_1_ca [3] $end
$var wire 1 c+ l1_1_ca [2] $end
$var wire 1 d+ l1_1_ca [1] $end
$var wire 1 e+ l1_1_ca [0] $end
$var wire 1 f+ l1_2_0 [39] $end
$var wire 1 g+ l1_2_0 [38] $end
$var wire 1 h+ l1_2_0 [37] $end
$var wire 1 i+ l1_2_0 [36] $end
$var wire 1 j+ l1_2_0 [35] $end
$var wire 1 k+ l1_2_0 [34] $end
$var wire 1 l+ l1_2_0 [33] $end
$var wire 1 m+ l1_2_0 [32] $end
$var wire 1 n+ l1_2_0 [31] $end
$var wire 1 o+ l1_2_0 [30] $end
$var wire 1 p+ l1_2_0 [29] $end
$var wire 1 q+ l1_2_0 [28] $end
$var wire 1 r+ l1_2_0 [27] $end
$var wire 1 s+ l1_2_0 [26] $end
$var wire 1 t+ l1_2_0 [25] $end
$var wire 1 u+ l1_2_0 [24] $end
$var wire 1 v+ l1_2_0 [23] $end
$var wire 1 w+ l1_2_0 [22] $end
$var wire 1 x+ l1_2_0 [21] $end
$var wire 1 y+ l1_2_0 [20] $end
$var wire 1 z+ l1_2_0 [19] $end
$var wire 1 {+ l1_2_0 [18] $end
$var wire 1 |+ l1_2_0 [17] $end
$var wire 1 }+ l1_2_0 [16] $end
$var wire 1 ~+ l1_2_0 [15] $end
$var wire 1 !, l1_2_0 [14] $end
$var wire 1 ", l1_2_0 [13] $end
$var wire 1 #, l1_2_0 [12] $end
$var wire 1 $, l1_2_0 [11] $end
$var wire 1 %, l1_2_0 [10] $end
$var wire 1 &, l1_2_0 [9] $end
$var wire 1 ', l1_2_0 [8] $end
$var wire 1 (, l1_2_0 [7] $end
$var wire 1 ), l1_2_0 [6] $end
$var wire 1 *, l1_2_0 [5] $end
$var wire 1 +, l1_2_0 [4] $end
$var wire 1 ,, l1_2_0 [3] $end
$var wire 1 -, l1_2_0 [2] $end
$var wire 1 ., l1_2_0 [1] $end
$var wire 1 /, l1_2_0 [0] $end
$var wire 1 0, l1_2_1 [39] $end
$var wire 1 1, l1_2_1 [38] $end
$var wire 1 2, l1_2_1 [37] $end
$var wire 1 3, l1_2_1 [36] $end
$var wire 1 4, l1_2_1 [35] $end
$var wire 1 5, l1_2_1 [34] $end
$var wire 1 6, l1_2_1 [33] $end
$var wire 1 7, l1_2_1 [32] $end
$var wire 1 8, l1_2_1 [31] $end
$var wire 1 9, l1_2_1 [30] $end
$var wire 1 :, l1_2_1 [29] $end
$var wire 1 ;, l1_2_1 [28] $end
$var wire 1 <, l1_2_1 [27] $end
$var wire 1 =, l1_2_1 [26] $end
$var wire 1 >, l1_2_1 [25] $end
$var wire 1 ?, l1_2_1 [24] $end
$var wire 1 @, l1_2_1 [23] $end
$var wire 1 A, l1_2_1 [22] $end
$var wire 1 B, l1_2_1 [21] $end
$var wire 1 C, l1_2_1 [20] $end
$var wire 1 D, l1_2_1 [19] $end
$var wire 1 E, l1_2_1 [18] $end
$var wire 1 F, l1_2_1 [17] $end
$var wire 1 G, l1_2_1 [16] $end
$var wire 1 H, l1_2_1 [15] $end
$var wire 1 I, l1_2_1 [14] $end
$var wire 1 J, l1_2_1 [13] $end
$var wire 1 K, l1_2_1 [12] $end
$var wire 1 L, l1_2_1 [11] $end
$var wire 1 M, l1_2_1 [10] $end
$var wire 1 N, l1_2_1 [9] $end
$var wire 1 O, l1_2_1 [8] $end
$var wire 1 P, l1_2_1 [7] $end
$var wire 1 Q, l1_2_1 [6] $end
$var wire 1 R, l1_2_1 [5] $end
$var wire 1 S, l1_2_1 [4] $end
$var wire 1 T, l1_2_1 [3] $end
$var wire 1 U, l1_2_1 [2] $end
$var wire 1 V, l1_2_1 [1] $end
$var wire 1 W, l1_2_1 [0] $end
$var wire 1 X, l1_2_2 [39] $end
$var wire 1 Y, l1_2_2 [38] $end
$var wire 1 Z, l1_2_2 [37] $end
$var wire 1 [, l1_2_2 [36] $end
$var wire 1 \, l1_2_2 [35] $end
$var wire 1 ], l1_2_2 [34] $end
$var wire 1 ^, l1_2_2 [33] $end
$var wire 1 _, l1_2_2 [32] $end
$var wire 1 `, l1_2_2 [31] $end
$var wire 1 a, l1_2_2 [30] $end
$var wire 1 b, l1_2_2 [29] $end
$var wire 1 c, l1_2_2 [28] $end
$var wire 1 d, l1_2_2 [27] $end
$var wire 1 e, l1_2_2 [26] $end
$var wire 1 f, l1_2_2 [25] $end
$var wire 1 g, l1_2_2 [24] $end
$var wire 1 h, l1_2_2 [23] $end
$var wire 1 i, l1_2_2 [22] $end
$var wire 1 j, l1_2_2 [21] $end
$var wire 1 k, l1_2_2 [20] $end
$var wire 1 l, l1_2_2 [19] $end
$var wire 1 m, l1_2_2 [18] $end
$var wire 1 n, l1_2_2 [17] $end
$var wire 1 o, l1_2_2 [16] $end
$var wire 1 p, l1_2_2 [15] $end
$var wire 1 q, l1_2_2 [14] $end
$var wire 1 r, l1_2_2 [13] $end
$var wire 1 s, l1_2_2 [12] $end
$var wire 1 t, l1_2_2 [11] $end
$var wire 1 u, l1_2_2 [10] $end
$var wire 1 v, l1_2_2 [9] $end
$var wire 1 w, l1_2_2 [8] $end
$var wire 1 x, l1_2_2 [7] $end
$var wire 1 y, l1_2_2 [6] $end
$var wire 1 z, l1_2_2 [5] $end
$var wire 1 {, l1_2_2 [4] $end
$var wire 1 |, l1_2_2 [3] $end
$var wire 1 }, l1_2_2 [2] $end
$var wire 1 ~, l1_2_2 [1] $end
$var wire 1 !- l1_2_2 [0] $end
$var wire 1 "- l1_2_cin [39] $end
$var wire 1 #- l1_2_cin [38] $end
$var wire 1 $- l1_2_cin [37] $end
$var wire 1 %- l1_2_cin [36] $end
$var wire 1 &- l1_2_cin [35] $end
$var wire 1 '- l1_2_cin [34] $end
$var wire 1 (- l1_2_cin [33] $end
$var wire 1 )- l1_2_cin [32] $end
$var wire 1 *- l1_2_cin [31] $end
$var wire 1 +- l1_2_cin [30] $end
$var wire 1 ,- l1_2_cin [29] $end
$var wire 1 -- l1_2_cin [28] $end
$var wire 1 .- l1_2_cin [27] $end
$var wire 1 /- l1_2_cin [26] $end
$var wire 1 0- l1_2_cin [25] $end
$var wire 1 1- l1_2_cin [24] $end
$var wire 1 2- l1_2_cin [23] $end
$var wire 1 3- l1_2_cin [22] $end
$var wire 1 4- l1_2_cin [21] $end
$var wire 1 5- l1_2_cin [20] $end
$var wire 1 6- l1_2_cin [19] $end
$var wire 1 7- l1_2_cin [18] $end
$var wire 1 8- l1_2_cin [17] $end
$var wire 1 9- l1_2_cin [16] $end
$var wire 1 :- l1_2_cin [15] $end
$var wire 1 ;- l1_2_cin [14] $end
$var wire 1 <- l1_2_cin [13] $end
$var wire 1 =- l1_2_cin [12] $end
$var wire 1 >- l1_2_cin [11] $end
$var wire 1 ?- l1_2_cin [10] $end
$var wire 1 @- l1_2_cin [9] $end
$var wire 1 A- l1_2_cin [8] $end
$var wire 1 B- l1_2_cin [7] $end
$var wire 1 C- l1_2_cin [6] $end
$var wire 1 D- l1_2_cin [5] $end
$var wire 1 E- l1_2_cin [4] $end
$var wire 1 F- l1_2_cin [3] $end
$var wire 1 G- l1_2_cin [2] $end
$var wire 1 H- l1_2_cin [1] $end
$var wire 1 I- l1_2_cin [0] $end
$var wire 1 J- l1_2_cout [39] $end
$var wire 1 K- l1_2_cout [38] $end
$var wire 1 L- l1_2_cout [37] $end
$var wire 1 M- l1_2_cout [36] $end
$var wire 1 N- l1_2_cout [35] $end
$var wire 1 O- l1_2_cout [34] $end
$var wire 1 P- l1_2_cout [33] $end
$var wire 1 Q- l1_2_cout [32] $end
$var wire 1 R- l1_2_cout [31] $end
$var wire 1 S- l1_2_cout [30] $end
$var wire 1 T- l1_2_cout [29] $end
$var wire 1 U- l1_2_cout [28] $end
$var wire 1 V- l1_2_cout [27] $end
$var wire 1 W- l1_2_cout [26] $end
$var wire 1 X- l1_2_cout [25] $end
$var wire 1 Y- l1_2_cout [24] $end
$var wire 1 Z- l1_2_cout [23] $end
$var wire 1 [- l1_2_cout [22] $end
$var wire 1 \- l1_2_cout [21] $end
$var wire 1 ]- l1_2_cout [20] $end
$var wire 1 ^- l1_2_cout [19] $end
$var wire 1 _- l1_2_cout [18] $end
$var wire 1 `- l1_2_cout [17] $end
$var wire 1 a- l1_2_cout [16] $end
$var wire 1 b- l1_2_cout [15] $end
$var wire 1 c- l1_2_cout [14] $end
$var wire 1 d- l1_2_cout [13] $end
$var wire 1 e- l1_2_cout [12] $end
$var wire 1 f- l1_2_cout [11] $end
$var wire 1 g- l1_2_cout [10] $end
$var wire 1 h- l1_2_cout [9] $end
$var wire 1 i- l1_2_cout [8] $end
$var wire 1 j- l1_2_cout [7] $end
$var wire 1 k- l1_2_cout [6] $end
$var wire 1 l- l1_2_cout [5] $end
$var wire 1 m- l1_2_cout [4] $end
$var wire 1 n- l1_2_cout [3] $end
$var wire 1 o- l1_2_cout [2] $end
$var wire 1 p- l1_2_cout [1] $end
$var wire 1 q- l1_2_cout [0] $end
$var wire 1 r- l1_2_s [39] $end
$var wire 1 s- l1_2_s [38] $end
$var wire 1 t- l1_2_s [37] $end
$var wire 1 u- l1_2_s [36] $end
$var wire 1 v- l1_2_s [35] $end
$var wire 1 w- l1_2_s [34] $end
$var wire 1 x- l1_2_s [33] $end
$var wire 1 y- l1_2_s [32] $end
$var wire 1 z- l1_2_s [31] $end
$var wire 1 {- l1_2_s [30] $end
$var wire 1 |- l1_2_s [29] $end
$var wire 1 }- l1_2_s [28] $end
$var wire 1 ~- l1_2_s [27] $end
$var wire 1 !. l1_2_s [26] $end
$var wire 1 ". l1_2_s [25] $end
$var wire 1 #. l1_2_s [24] $end
$var wire 1 $. l1_2_s [23] $end
$var wire 1 %. l1_2_s [22] $end
$var wire 1 &. l1_2_s [21] $end
$var wire 1 '. l1_2_s [20] $end
$var wire 1 (. l1_2_s [19] $end
$var wire 1 ). l1_2_s [18] $end
$var wire 1 *. l1_2_s [17] $end
$var wire 1 +. l1_2_s [16] $end
$var wire 1 ,. l1_2_s [15] $end
$var wire 1 -. l1_2_s [14] $end
$var wire 1 .. l1_2_s [13] $end
$var wire 1 /. l1_2_s [12] $end
$var wire 1 0. l1_2_s [11] $end
$var wire 1 1. l1_2_s [10] $end
$var wire 1 2. l1_2_s [9] $end
$var wire 1 3. l1_2_s [8] $end
$var wire 1 4. l1_2_s [7] $end
$var wire 1 5. l1_2_s [6] $end
$var wire 1 6. l1_2_s [5] $end
$var wire 1 7. l1_2_s [4] $end
$var wire 1 8. l1_2_s [3] $end
$var wire 1 9. l1_2_s [2] $end
$var wire 1 :. l1_2_s [1] $end
$var wire 1 ;. l1_2_s [0] $end
$var wire 1 <. l1_2_ca [39] $end
$var wire 1 =. l1_2_ca [38] $end
$var wire 1 >. l1_2_ca [37] $end
$var wire 1 ?. l1_2_ca [36] $end
$var wire 1 @. l1_2_ca [35] $end
$var wire 1 A. l1_2_ca [34] $end
$var wire 1 B. l1_2_ca [33] $end
$var wire 1 C. l1_2_ca [32] $end
$var wire 1 D. l1_2_ca [31] $end
$var wire 1 E. l1_2_ca [30] $end
$var wire 1 F. l1_2_ca [29] $end
$var wire 1 G. l1_2_ca [28] $end
$var wire 1 H. l1_2_ca [27] $end
$var wire 1 I. l1_2_ca [26] $end
$var wire 1 J. l1_2_ca [25] $end
$var wire 1 K. l1_2_ca [24] $end
$var wire 1 L. l1_2_ca [23] $end
$var wire 1 M. l1_2_ca [22] $end
$var wire 1 N. l1_2_ca [21] $end
$var wire 1 O. l1_2_ca [20] $end
$var wire 1 P. l1_2_ca [19] $end
$var wire 1 Q. l1_2_ca [18] $end
$var wire 1 R. l1_2_ca [17] $end
$var wire 1 S. l1_2_ca [16] $end
$var wire 1 T. l1_2_ca [15] $end
$var wire 1 U. l1_2_ca [14] $end
$var wire 1 V. l1_2_ca [13] $end
$var wire 1 W. l1_2_ca [12] $end
$var wire 1 X. l1_2_ca [11] $end
$var wire 1 Y. l1_2_ca [10] $end
$var wire 1 Z. l1_2_ca [9] $end
$var wire 1 [. l1_2_ca [8] $end
$var wire 1 \. l1_2_ca [7] $end
$var wire 1 ]. l1_2_ca [6] $end
$var wire 1 ^. l1_2_ca [5] $end
$var wire 1 _. l1_2_ca [4] $end
$var wire 1 `. l1_2_ca [3] $end
$var wire 1 a. l1_2_ca [2] $end
$var wire 1 b. l1_2_ca [1] $end
$var wire 1 c. l1_2_ca [0] $end
$var wire 1 d. l1_3_0 [39] $end
$var wire 1 e. l1_3_0 [38] $end
$var wire 1 f. l1_3_0 [37] $end
$var wire 1 g. l1_3_0 [36] $end
$var wire 1 h. l1_3_0 [35] $end
$var wire 1 i. l1_3_0 [34] $end
$var wire 1 j. l1_3_0 [33] $end
$var wire 1 k. l1_3_0 [32] $end
$var wire 1 l. l1_3_0 [31] $end
$var wire 1 m. l1_3_0 [30] $end
$var wire 1 n. l1_3_0 [29] $end
$var wire 1 o. l1_3_0 [28] $end
$var wire 1 p. l1_3_0 [27] $end
$var wire 1 q. l1_3_0 [26] $end
$var wire 1 r. l1_3_0 [25] $end
$var wire 1 s. l1_3_0 [24] $end
$var wire 1 t. l1_3_0 [23] $end
$var wire 1 u. l1_3_0 [22] $end
$var wire 1 v. l1_3_0 [21] $end
$var wire 1 w. l1_3_0 [20] $end
$var wire 1 x. l1_3_0 [19] $end
$var wire 1 y. l1_3_0 [18] $end
$var wire 1 z. l1_3_0 [17] $end
$var wire 1 {. l1_3_0 [16] $end
$var wire 1 |. l1_3_0 [15] $end
$var wire 1 }. l1_3_0 [14] $end
$var wire 1 ~. l1_3_0 [13] $end
$var wire 1 !/ l1_3_0 [12] $end
$var wire 1 "/ l1_3_0 [11] $end
$var wire 1 #/ l1_3_0 [10] $end
$var wire 1 $/ l1_3_0 [9] $end
$var wire 1 %/ l1_3_0 [8] $end
$var wire 1 &/ l1_3_0 [7] $end
$var wire 1 '/ l1_3_0 [6] $end
$var wire 1 (/ l1_3_0 [5] $end
$var wire 1 )/ l1_3_0 [4] $end
$var wire 1 */ l1_3_0 [3] $end
$var wire 1 +/ l1_3_0 [2] $end
$var wire 1 ,/ l1_3_0 [1] $end
$var wire 1 -/ l1_3_0 [0] $end
$var wire 1 ./ l1_3_1 [39] $end
$var wire 1 // l1_3_1 [38] $end
$var wire 1 0/ l1_3_1 [37] $end
$var wire 1 1/ l1_3_1 [36] $end
$var wire 1 2/ l1_3_1 [35] $end
$var wire 1 3/ l1_3_1 [34] $end
$var wire 1 4/ l1_3_1 [33] $end
$var wire 1 5/ l1_3_1 [32] $end
$var wire 1 6/ l1_3_1 [31] $end
$var wire 1 7/ l1_3_1 [30] $end
$var wire 1 8/ l1_3_1 [29] $end
$var wire 1 9/ l1_3_1 [28] $end
$var wire 1 :/ l1_3_1 [27] $end
$var wire 1 ;/ l1_3_1 [26] $end
$var wire 1 </ l1_3_1 [25] $end
$var wire 1 =/ l1_3_1 [24] $end
$var wire 1 >/ l1_3_1 [23] $end
$var wire 1 ?/ l1_3_1 [22] $end
$var wire 1 @/ l1_3_1 [21] $end
$var wire 1 A/ l1_3_1 [20] $end
$var wire 1 B/ l1_3_1 [19] $end
$var wire 1 C/ l1_3_1 [18] $end
$var wire 1 D/ l1_3_1 [17] $end
$var wire 1 E/ l1_3_1 [16] $end
$var wire 1 F/ l1_3_1 [15] $end
$var wire 1 G/ l1_3_1 [14] $end
$var wire 1 H/ l1_3_1 [13] $end
$var wire 1 I/ l1_3_1 [12] $end
$var wire 1 J/ l1_3_1 [11] $end
$var wire 1 K/ l1_3_1 [10] $end
$var wire 1 L/ l1_3_1 [9] $end
$var wire 1 M/ l1_3_1 [8] $end
$var wire 1 N/ l1_3_1 [7] $end
$var wire 1 O/ l1_3_1 [6] $end
$var wire 1 P/ l1_3_1 [5] $end
$var wire 1 Q/ l1_3_1 [4] $end
$var wire 1 R/ l1_3_1 [3] $end
$var wire 1 S/ l1_3_1 [2] $end
$var wire 1 T/ l1_3_1 [1] $end
$var wire 1 U/ l1_3_1 [0] $end
$var wire 1 V/ l1_3_2 [39] $end
$var wire 1 W/ l1_3_2 [38] $end
$var wire 1 X/ l1_3_2 [37] $end
$var wire 1 Y/ l1_3_2 [36] $end
$var wire 1 Z/ l1_3_2 [35] $end
$var wire 1 [/ l1_3_2 [34] $end
$var wire 1 \/ l1_3_2 [33] $end
$var wire 1 ]/ l1_3_2 [32] $end
$var wire 1 ^/ l1_3_2 [31] $end
$var wire 1 _/ l1_3_2 [30] $end
$var wire 1 `/ l1_3_2 [29] $end
$var wire 1 a/ l1_3_2 [28] $end
$var wire 1 b/ l1_3_2 [27] $end
$var wire 1 c/ l1_3_2 [26] $end
$var wire 1 d/ l1_3_2 [25] $end
$var wire 1 e/ l1_3_2 [24] $end
$var wire 1 f/ l1_3_2 [23] $end
$var wire 1 g/ l1_3_2 [22] $end
$var wire 1 h/ l1_3_2 [21] $end
$var wire 1 i/ l1_3_2 [20] $end
$var wire 1 j/ l1_3_2 [19] $end
$var wire 1 k/ l1_3_2 [18] $end
$var wire 1 l/ l1_3_2 [17] $end
$var wire 1 m/ l1_3_2 [16] $end
$var wire 1 n/ l1_3_2 [15] $end
$var wire 1 o/ l1_3_2 [14] $end
$var wire 1 p/ l1_3_2 [13] $end
$var wire 1 q/ l1_3_2 [12] $end
$var wire 1 r/ l1_3_2 [11] $end
$var wire 1 s/ l1_3_2 [10] $end
$var wire 1 t/ l1_3_2 [9] $end
$var wire 1 u/ l1_3_2 [8] $end
$var wire 1 v/ l1_3_2 [7] $end
$var wire 1 w/ l1_3_2 [6] $end
$var wire 1 x/ l1_3_2 [5] $end
$var wire 1 y/ l1_3_2 [4] $end
$var wire 1 z/ l1_3_2 [3] $end
$var wire 1 {/ l1_3_2 [2] $end
$var wire 1 |/ l1_3_2 [1] $end
$var wire 1 }/ l1_3_2 [0] $end
$var wire 1 ~/ l1_3_cin [39] $end
$var wire 1 !0 l1_3_cin [38] $end
$var wire 1 "0 l1_3_cin [37] $end
$var wire 1 #0 l1_3_cin [36] $end
$var wire 1 $0 l1_3_cin [35] $end
$var wire 1 %0 l1_3_cin [34] $end
$var wire 1 &0 l1_3_cin [33] $end
$var wire 1 '0 l1_3_cin [32] $end
$var wire 1 (0 l1_3_cin [31] $end
$var wire 1 )0 l1_3_cin [30] $end
$var wire 1 *0 l1_3_cin [29] $end
$var wire 1 +0 l1_3_cin [28] $end
$var wire 1 ,0 l1_3_cin [27] $end
$var wire 1 -0 l1_3_cin [26] $end
$var wire 1 .0 l1_3_cin [25] $end
$var wire 1 /0 l1_3_cin [24] $end
$var wire 1 00 l1_3_cin [23] $end
$var wire 1 10 l1_3_cin [22] $end
$var wire 1 20 l1_3_cin [21] $end
$var wire 1 30 l1_3_cin [20] $end
$var wire 1 40 l1_3_cin [19] $end
$var wire 1 50 l1_3_cin [18] $end
$var wire 1 60 l1_3_cin [17] $end
$var wire 1 70 l1_3_cin [16] $end
$var wire 1 80 l1_3_cin [15] $end
$var wire 1 90 l1_3_cin [14] $end
$var wire 1 :0 l1_3_cin [13] $end
$var wire 1 ;0 l1_3_cin [12] $end
$var wire 1 <0 l1_3_cin [11] $end
$var wire 1 =0 l1_3_cin [10] $end
$var wire 1 >0 l1_3_cin [9] $end
$var wire 1 ?0 l1_3_cin [8] $end
$var wire 1 @0 l1_3_cin [7] $end
$var wire 1 A0 l1_3_cin [6] $end
$var wire 1 B0 l1_3_cin [5] $end
$var wire 1 C0 l1_3_cin [4] $end
$var wire 1 D0 l1_3_cin [3] $end
$var wire 1 E0 l1_3_cin [2] $end
$var wire 1 F0 l1_3_cin [1] $end
$var wire 1 G0 l1_3_cin [0] $end
$var wire 1 H0 l1_3_cout [39] $end
$var wire 1 I0 l1_3_cout [38] $end
$var wire 1 J0 l1_3_cout [37] $end
$var wire 1 K0 l1_3_cout [36] $end
$var wire 1 L0 l1_3_cout [35] $end
$var wire 1 M0 l1_3_cout [34] $end
$var wire 1 N0 l1_3_cout [33] $end
$var wire 1 O0 l1_3_cout [32] $end
$var wire 1 P0 l1_3_cout [31] $end
$var wire 1 Q0 l1_3_cout [30] $end
$var wire 1 R0 l1_3_cout [29] $end
$var wire 1 S0 l1_3_cout [28] $end
$var wire 1 T0 l1_3_cout [27] $end
$var wire 1 U0 l1_3_cout [26] $end
$var wire 1 V0 l1_3_cout [25] $end
$var wire 1 W0 l1_3_cout [24] $end
$var wire 1 X0 l1_3_cout [23] $end
$var wire 1 Y0 l1_3_cout [22] $end
$var wire 1 Z0 l1_3_cout [21] $end
$var wire 1 [0 l1_3_cout [20] $end
$var wire 1 \0 l1_3_cout [19] $end
$var wire 1 ]0 l1_3_cout [18] $end
$var wire 1 ^0 l1_3_cout [17] $end
$var wire 1 _0 l1_3_cout [16] $end
$var wire 1 `0 l1_3_cout [15] $end
$var wire 1 a0 l1_3_cout [14] $end
$var wire 1 b0 l1_3_cout [13] $end
$var wire 1 c0 l1_3_cout [12] $end
$var wire 1 d0 l1_3_cout [11] $end
$var wire 1 e0 l1_3_cout [10] $end
$var wire 1 f0 l1_3_cout [9] $end
$var wire 1 g0 l1_3_cout [8] $end
$var wire 1 h0 l1_3_cout [7] $end
$var wire 1 i0 l1_3_cout [6] $end
$var wire 1 j0 l1_3_cout [5] $end
$var wire 1 k0 l1_3_cout [4] $end
$var wire 1 l0 l1_3_cout [3] $end
$var wire 1 m0 l1_3_cout [2] $end
$var wire 1 n0 l1_3_cout [1] $end
$var wire 1 o0 l1_3_cout [0] $end
$var wire 1 p0 l1_3_s [39] $end
$var wire 1 q0 l1_3_s [38] $end
$var wire 1 r0 l1_3_s [37] $end
$var wire 1 s0 l1_3_s [36] $end
$var wire 1 t0 l1_3_s [35] $end
$var wire 1 u0 l1_3_s [34] $end
$var wire 1 v0 l1_3_s [33] $end
$var wire 1 w0 l1_3_s [32] $end
$var wire 1 x0 l1_3_s [31] $end
$var wire 1 y0 l1_3_s [30] $end
$var wire 1 z0 l1_3_s [29] $end
$var wire 1 {0 l1_3_s [28] $end
$var wire 1 |0 l1_3_s [27] $end
$var wire 1 }0 l1_3_s [26] $end
$var wire 1 ~0 l1_3_s [25] $end
$var wire 1 !1 l1_3_s [24] $end
$var wire 1 "1 l1_3_s [23] $end
$var wire 1 #1 l1_3_s [22] $end
$var wire 1 $1 l1_3_s [21] $end
$var wire 1 %1 l1_3_s [20] $end
$var wire 1 &1 l1_3_s [19] $end
$var wire 1 '1 l1_3_s [18] $end
$var wire 1 (1 l1_3_s [17] $end
$var wire 1 )1 l1_3_s [16] $end
$var wire 1 *1 l1_3_s [15] $end
$var wire 1 +1 l1_3_s [14] $end
$var wire 1 ,1 l1_3_s [13] $end
$var wire 1 -1 l1_3_s [12] $end
$var wire 1 .1 l1_3_s [11] $end
$var wire 1 /1 l1_3_s [10] $end
$var wire 1 01 l1_3_s [9] $end
$var wire 1 11 l1_3_s [8] $end
$var wire 1 21 l1_3_s [7] $end
$var wire 1 31 l1_3_s [6] $end
$var wire 1 41 l1_3_s [5] $end
$var wire 1 51 l1_3_s [4] $end
$var wire 1 61 l1_3_s [3] $end
$var wire 1 71 l1_3_s [2] $end
$var wire 1 81 l1_3_s [1] $end
$var wire 1 91 l1_3_s [0] $end
$var wire 1 :1 l1_3_ca [39] $end
$var wire 1 ;1 l1_3_ca [38] $end
$var wire 1 <1 l1_3_ca [37] $end
$var wire 1 =1 l1_3_ca [36] $end
$var wire 1 >1 l1_3_ca [35] $end
$var wire 1 ?1 l1_3_ca [34] $end
$var wire 1 @1 l1_3_ca [33] $end
$var wire 1 A1 l1_3_ca [32] $end
$var wire 1 B1 l1_3_ca [31] $end
$var wire 1 C1 l1_3_ca [30] $end
$var wire 1 D1 l1_3_ca [29] $end
$var wire 1 E1 l1_3_ca [28] $end
$var wire 1 F1 l1_3_ca [27] $end
$var wire 1 G1 l1_3_ca [26] $end
$var wire 1 H1 l1_3_ca [25] $end
$var wire 1 I1 l1_3_ca [24] $end
$var wire 1 J1 l1_3_ca [23] $end
$var wire 1 K1 l1_3_ca [22] $end
$var wire 1 L1 l1_3_ca [21] $end
$var wire 1 M1 l1_3_ca [20] $end
$var wire 1 N1 l1_3_ca [19] $end
$var wire 1 O1 l1_3_ca [18] $end
$var wire 1 P1 l1_3_ca [17] $end
$var wire 1 Q1 l1_3_ca [16] $end
$var wire 1 R1 l1_3_ca [15] $end
$var wire 1 S1 l1_3_ca [14] $end
$var wire 1 T1 l1_3_ca [13] $end
$var wire 1 U1 l1_3_ca [12] $end
$var wire 1 V1 l1_3_ca [11] $end
$var wire 1 W1 l1_3_ca [10] $end
$var wire 1 X1 l1_3_ca [9] $end
$var wire 1 Y1 l1_3_ca [8] $end
$var wire 1 Z1 l1_3_ca [7] $end
$var wire 1 [1 l1_3_ca [6] $end
$var wire 1 \1 l1_3_ca [5] $end
$var wire 1 ]1 l1_3_ca [4] $end
$var wire 1 ^1 l1_3_ca [3] $end
$var wire 1 _1 l1_3_ca [2] $end
$var wire 1 `1 l1_3_ca [1] $end
$var wire 1 a1 l1_3_ca [0] $end
$var wire 1 b1 l1_4_0 [39] $end
$var wire 1 c1 l1_4_0 [38] $end
$var wire 1 d1 l1_4_0 [37] $end
$var wire 1 e1 l1_4_0 [36] $end
$var wire 1 f1 l1_4_0 [35] $end
$var wire 1 g1 l1_4_0 [34] $end
$var wire 1 h1 l1_4_0 [33] $end
$var wire 1 i1 l1_4_0 [32] $end
$var wire 1 j1 l1_4_0 [31] $end
$var wire 1 k1 l1_4_0 [30] $end
$var wire 1 l1 l1_4_0 [29] $end
$var wire 1 m1 l1_4_0 [28] $end
$var wire 1 n1 l1_4_0 [27] $end
$var wire 1 o1 l1_4_0 [26] $end
$var wire 1 p1 l1_4_0 [25] $end
$var wire 1 q1 l1_4_0 [24] $end
$var wire 1 r1 l1_4_0 [23] $end
$var wire 1 s1 l1_4_0 [22] $end
$var wire 1 t1 l1_4_0 [21] $end
$var wire 1 u1 l1_4_0 [20] $end
$var wire 1 v1 l1_4_0 [19] $end
$var wire 1 w1 l1_4_0 [18] $end
$var wire 1 x1 l1_4_0 [17] $end
$var wire 1 y1 l1_4_0 [16] $end
$var wire 1 z1 l1_4_0 [15] $end
$var wire 1 {1 l1_4_0 [14] $end
$var wire 1 |1 l1_4_0 [13] $end
$var wire 1 }1 l1_4_0 [12] $end
$var wire 1 ~1 l1_4_0 [11] $end
$var wire 1 !2 l1_4_0 [10] $end
$var wire 1 "2 l1_4_0 [9] $end
$var wire 1 #2 l1_4_0 [8] $end
$var wire 1 $2 l1_4_0 [7] $end
$var wire 1 %2 l1_4_0 [6] $end
$var wire 1 &2 l1_4_0 [5] $end
$var wire 1 '2 l1_4_0 [4] $end
$var wire 1 (2 l1_4_0 [3] $end
$var wire 1 )2 l1_4_0 [2] $end
$var wire 1 *2 l1_4_0 [1] $end
$var wire 1 +2 l1_4_0 [0] $end
$var wire 1 ,2 l1_4_1 [39] $end
$var wire 1 -2 l1_4_1 [38] $end
$var wire 1 .2 l1_4_1 [37] $end
$var wire 1 /2 l1_4_1 [36] $end
$var wire 1 02 l1_4_1 [35] $end
$var wire 1 12 l1_4_1 [34] $end
$var wire 1 22 l1_4_1 [33] $end
$var wire 1 32 l1_4_1 [32] $end
$var wire 1 42 l1_4_1 [31] $end
$var wire 1 52 l1_4_1 [30] $end
$var wire 1 62 l1_4_1 [29] $end
$var wire 1 72 l1_4_1 [28] $end
$var wire 1 82 l1_4_1 [27] $end
$var wire 1 92 l1_4_1 [26] $end
$var wire 1 :2 l1_4_1 [25] $end
$var wire 1 ;2 l1_4_1 [24] $end
$var wire 1 <2 l1_4_1 [23] $end
$var wire 1 =2 l1_4_1 [22] $end
$var wire 1 >2 l1_4_1 [21] $end
$var wire 1 ?2 l1_4_1 [20] $end
$var wire 1 @2 l1_4_1 [19] $end
$var wire 1 A2 l1_4_1 [18] $end
$var wire 1 B2 l1_4_1 [17] $end
$var wire 1 C2 l1_4_1 [16] $end
$var wire 1 D2 l1_4_1 [15] $end
$var wire 1 E2 l1_4_1 [14] $end
$var wire 1 F2 l1_4_1 [13] $end
$var wire 1 G2 l1_4_1 [12] $end
$var wire 1 H2 l1_4_1 [11] $end
$var wire 1 I2 l1_4_1 [10] $end
$var wire 1 J2 l1_4_1 [9] $end
$var wire 1 K2 l1_4_1 [8] $end
$var wire 1 L2 l1_4_1 [7] $end
$var wire 1 M2 l1_4_1 [6] $end
$var wire 1 N2 l1_4_1 [5] $end
$var wire 1 O2 l1_4_1 [4] $end
$var wire 1 P2 l1_4_1 [3] $end
$var wire 1 Q2 l1_4_1 [2] $end
$var wire 1 R2 l1_4_1 [1] $end
$var wire 1 S2 l1_4_1 [0] $end
$var wire 1 T2 l1_4_2 [39] $end
$var wire 1 U2 l1_4_2 [38] $end
$var wire 1 V2 l1_4_2 [37] $end
$var wire 1 W2 l1_4_2 [36] $end
$var wire 1 X2 l1_4_2 [35] $end
$var wire 1 Y2 l1_4_2 [34] $end
$var wire 1 Z2 l1_4_2 [33] $end
$var wire 1 [2 l1_4_2 [32] $end
$var wire 1 \2 l1_4_2 [31] $end
$var wire 1 ]2 l1_4_2 [30] $end
$var wire 1 ^2 l1_4_2 [29] $end
$var wire 1 _2 l1_4_2 [28] $end
$var wire 1 `2 l1_4_2 [27] $end
$var wire 1 a2 l1_4_2 [26] $end
$var wire 1 b2 l1_4_2 [25] $end
$var wire 1 c2 l1_4_2 [24] $end
$var wire 1 d2 l1_4_2 [23] $end
$var wire 1 e2 l1_4_2 [22] $end
$var wire 1 f2 l1_4_2 [21] $end
$var wire 1 g2 l1_4_2 [20] $end
$var wire 1 h2 l1_4_2 [19] $end
$var wire 1 i2 l1_4_2 [18] $end
$var wire 1 j2 l1_4_2 [17] $end
$var wire 1 k2 l1_4_2 [16] $end
$var wire 1 l2 l1_4_2 [15] $end
$var wire 1 m2 l1_4_2 [14] $end
$var wire 1 n2 l1_4_2 [13] $end
$var wire 1 o2 l1_4_2 [12] $end
$var wire 1 p2 l1_4_2 [11] $end
$var wire 1 q2 l1_4_2 [10] $end
$var wire 1 r2 l1_4_2 [9] $end
$var wire 1 s2 l1_4_2 [8] $end
$var wire 1 t2 l1_4_2 [7] $end
$var wire 1 u2 l1_4_2 [6] $end
$var wire 1 v2 l1_4_2 [5] $end
$var wire 1 w2 l1_4_2 [4] $end
$var wire 1 x2 l1_4_2 [3] $end
$var wire 1 y2 l1_4_2 [2] $end
$var wire 1 z2 l1_4_2 [1] $end
$var wire 1 {2 l1_4_2 [0] $end
$var wire 1 |2 l1_4_cin [39] $end
$var wire 1 }2 l1_4_cin [38] $end
$var wire 1 ~2 l1_4_cin [37] $end
$var wire 1 !3 l1_4_cin [36] $end
$var wire 1 "3 l1_4_cin [35] $end
$var wire 1 #3 l1_4_cin [34] $end
$var wire 1 $3 l1_4_cin [33] $end
$var wire 1 %3 l1_4_cin [32] $end
$var wire 1 &3 l1_4_cin [31] $end
$var wire 1 '3 l1_4_cin [30] $end
$var wire 1 (3 l1_4_cin [29] $end
$var wire 1 )3 l1_4_cin [28] $end
$var wire 1 *3 l1_4_cin [27] $end
$var wire 1 +3 l1_4_cin [26] $end
$var wire 1 ,3 l1_4_cin [25] $end
$var wire 1 -3 l1_4_cin [24] $end
$var wire 1 .3 l1_4_cin [23] $end
$var wire 1 /3 l1_4_cin [22] $end
$var wire 1 03 l1_4_cin [21] $end
$var wire 1 13 l1_4_cin [20] $end
$var wire 1 23 l1_4_cin [19] $end
$var wire 1 33 l1_4_cin [18] $end
$var wire 1 43 l1_4_cin [17] $end
$var wire 1 53 l1_4_cin [16] $end
$var wire 1 63 l1_4_cin [15] $end
$var wire 1 73 l1_4_cin [14] $end
$var wire 1 83 l1_4_cin [13] $end
$var wire 1 93 l1_4_cin [12] $end
$var wire 1 :3 l1_4_cin [11] $end
$var wire 1 ;3 l1_4_cin [10] $end
$var wire 1 <3 l1_4_cin [9] $end
$var wire 1 =3 l1_4_cin [8] $end
$var wire 1 >3 l1_4_cin [7] $end
$var wire 1 ?3 l1_4_cin [6] $end
$var wire 1 @3 l1_4_cin [5] $end
$var wire 1 A3 l1_4_cin [4] $end
$var wire 1 B3 l1_4_cin [3] $end
$var wire 1 C3 l1_4_cin [2] $end
$var wire 1 D3 l1_4_cin [1] $end
$var wire 1 E3 l1_4_cin [0] $end
$var wire 1 F3 l1_4_cout [39] $end
$var wire 1 G3 l1_4_cout [38] $end
$var wire 1 H3 l1_4_cout [37] $end
$var wire 1 I3 l1_4_cout [36] $end
$var wire 1 J3 l1_4_cout [35] $end
$var wire 1 K3 l1_4_cout [34] $end
$var wire 1 L3 l1_4_cout [33] $end
$var wire 1 M3 l1_4_cout [32] $end
$var wire 1 N3 l1_4_cout [31] $end
$var wire 1 O3 l1_4_cout [30] $end
$var wire 1 P3 l1_4_cout [29] $end
$var wire 1 Q3 l1_4_cout [28] $end
$var wire 1 R3 l1_4_cout [27] $end
$var wire 1 S3 l1_4_cout [26] $end
$var wire 1 T3 l1_4_cout [25] $end
$var wire 1 U3 l1_4_cout [24] $end
$var wire 1 V3 l1_4_cout [23] $end
$var wire 1 W3 l1_4_cout [22] $end
$var wire 1 X3 l1_4_cout [21] $end
$var wire 1 Y3 l1_4_cout [20] $end
$var wire 1 Z3 l1_4_cout [19] $end
$var wire 1 [3 l1_4_cout [18] $end
$var wire 1 \3 l1_4_cout [17] $end
$var wire 1 ]3 l1_4_cout [16] $end
$var wire 1 ^3 l1_4_cout [15] $end
$var wire 1 _3 l1_4_cout [14] $end
$var wire 1 `3 l1_4_cout [13] $end
$var wire 1 a3 l1_4_cout [12] $end
$var wire 1 b3 l1_4_cout [11] $end
$var wire 1 c3 l1_4_cout [10] $end
$var wire 1 d3 l1_4_cout [9] $end
$var wire 1 e3 l1_4_cout [8] $end
$var wire 1 f3 l1_4_cout [7] $end
$var wire 1 g3 l1_4_cout [6] $end
$var wire 1 h3 l1_4_cout [5] $end
$var wire 1 i3 l1_4_cout [4] $end
$var wire 1 j3 l1_4_cout [3] $end
$var wire 1 k3 l1_4_cout [2] $end
$var wire 1 l3 l1_4_cout [1] $end
$var wire 1 m3 l1_4_cout [0] $end
$var wire 1 n3 l1_4_s [39] $end
$var wire 1 o3 l1_4_s [38] $end
$var wire 1 p3 l1_4_s [37] $end
$var wire 1 q3 l1_4_s [36] $end
$var wire 1 r3 l1_4_s [35] $end
$var wire 1 s3 l1_4_s [34] $end
$var wire 1 t3 l1_4_s [33] $end
$var wire 1 u3 l1_4_s [32] $end
$var wire 1 v3 l1_4_s [31] $end
$var wire 1 w3 l1_4_s [30] $end
$var wire 1 x3 l1_4_s [29] $end
$var wire 1 y3 l1_4_s [28] $end
$var wire 1 z3 l1_4_s [27] $end
$var wire 1 {3 l1_4_s [26] $end
$var wire 1 |3 l1_4_s [25] $end
$var wire 1 }3 l1_4_s [24] $end
$var wire 1 ~3 l1_4_s [23] $end
$var wire 1 !4 l1_4_s [22] $end
$var wire 1 "4 l1_4_s [21] $end
$var wire 1 #4 l1_4_s [20] $end
$var wire 1 $4 l1_4_s [19] $end
$var wire 1 %4 l1_4_s [18] $end
$var wire 1 &4 l1_4_s [17] $end
$var wire 1 '4 l1_4_s [16] $end
$var wire 1 (4 l1_4_s [15] $end
$var wire 1 )4 l1_4_s [14] $end
$var wire 1 *4 l1_4_s [13] $end
$var wire 1 +4 l1_4_s [12] $end
$var wire 1 ,4 l1_4_s [11] $end
$var wire 1 -4 l1_4_s [10] $end
$var wire 1 .4 l1_4_s [9] $end
$var wire 1 /4 l1_4_s [8] $end
$var wire 1 04 l1_4_s [7] $end
$var wire 1 14 l1_4_s [6] $end
$var wire 1 24 l1_4_s [5] $end
$var wire 1 34 l1_4_s [4] $end
$var wire 1 44 l1_4_s [3] $end
$var wire 1 54 l1_4_s [2] $end
$var wire 1 64 l1_4_s [1] $end
$var wire 1 74 l1_4_s [0] $end
$var wire 1 84 l1_4_ca [39] $end
$var wire 1 94 l1_4_ca [38] $end
$var wire 1 :4 l1_4_ca [37] $end
$var wire 1 ;4 l1_4_ca [36] $end
$var wire 1 <4 l1_4_ca [35] $end
$var wire 1 =4 l1_4_ca [34] $end
$var wire 1 >4 l1_4_ca [33] $end
$var wire 1 ?4 l1_4_ca [32] $end
$var wire 1 @4 l1_4_ca [31] $end
$var wire 1 A4 l1_4_ca [30] $end
$var wire 1 B4 l1_4_ca [29] $end
$var wire 1 C4 l1_4_ca [28] $end
$var wire 1 D4 l1_4_ca [27] $end
$var wire 1 E4 l1_4_ca [26] $end
$var wire 1 F4 l1_4_ca [25] $end
$var wire 1 G4 l1_4_ca [24] $end
$var wire 1 H4 l1_4_ca [23] $end
$var wire 1 I4 l1_4_ca [22] $end
$var wire 1 J4 l1_4_ca [21] $end
$var wire 1 K4 l1_4_ca [20] $end
$var wire 1 L4 l1_4_ca [19] $end
$var wire 1 M4 l1_4_ca [18] $end
$var wire 1 N4 l1_4_ca [17] $end
$var wire 1 O4 l1_4_ca [16] $end
$var wire 1 P4 l1_4_ca [15] $end
$var wire 1 Q4 l1_4_ca [14] $end
$var wire 1 R4 l1_4_ca [13] $end
$var wire 1 S4 l1_4_ca [12] $end
$var wire 1 T4 l1_4_ca [11] $end
$var wire 1 U4 l1_4_ca [10] $end
$var wire 1 V4 l1_4_ca [9] $end
$var wire 1 W4 l1_4_ca [8] $end
$var wire 1 X4 l1_4_ca [7] $end
$var wire 1 Y4 l1_4_ca [6] $end
$var wire 1 Z4 l1_4_ca [5] $end
$var wire 1 [4 l1_4_ca [4] $end
$var wire 1 \4 l1_4_ca [3] $end
$var wire 1 ]4 l1_4_ca [2] $end
$var wire 1 ^4 l1_4_ca [1] $end
$var wire 1 _4 l1_4_ca [0] $end
$var wire 1 `4 l1_5_0 [39] $end
$var wire 1 a4 l1_5_0 [38] $end
$var wire 1 b4 l1_5_0 [37] $end
$var wire 1 c4 l1_5_0 [36] $end
$var wire 1 d4 l1_5_0 [35] $end
$var wire 1 e4 l1_5_0 [34] $end
$var wire 1 f4 l1_5_0 [33] $end
$var wire 1 g4 l1_5_0 [32] $end
$var wire 1 h4 l1_5_0 [31] $end
$var wire 1 i4 l1_5_0 [30] $end
$var wire 1 j4 l1_5_0 [29] $end
$var wire 1 k4 l1_5_0 [28] $end
$var wire 1 l4 l1_5_0 [27] $end
$var wire 1 m4 l1_5_0 [26] $end
$var wire 1 n4 l1_5_0 [25] $end
$var wire 1 o4 l1_5_0 [24] $end
$var wire 1 p4 l1_5_0 [23] $end
$var wire 1 q4 l1_5_0 [22] $end
$var wire 1 r4 l1_5_0 [21] $end
$var wire 1 s4 l1_5_0 [20] $end
$var wire 1 t4 l1_5_0 [19] $end
$var wire 1 u4 l1_5_0 [18] $end
$var wire 1 v4 l1_5_0 [17] $end
$var wire 1 w4 l1_5_0 [16] $end
$var wire 1 x4 l1_5_0 [15] $end
$var wire 1 y4 l1_5_0 [14] $end
$var wire 1 z4 l1_5_0 [13] $end
$var wire 1 {4 l1_5_0 [12] $end
$var wire 1 |4 l1_5_0 [11] $end
$var wire 1 }4 l1_5_0 [10] $end
$var wire 1 ~4 l1_5_0 [9] $end
$var wire 1 !5 l1_5_0 [8] $end
$var wire 1 "5 l1_5_0 [7] $end
$var wire 1 #5 l1_5_0 [6] $end
$var wire 1 $5 l1_5_0 [5] $end
$var wire 1 %5 l1_5_0 [4] $end
$var wire 1 &5 l1_5_0 [3] $end
$var wire 1 '5 l1_5_0 [2] $end
$var wire 1 (5 l1_5_0 [1] $end
$var wire 1 )5 l1_5_0 [0] $end
$var wire 1 *5 l1_5_1 [39] $end
$var wire 1 +5 l1_5_1 [38] $end
$var wire 1 ,5 l1_5_1 [37] $end
$var wire 1 -5 l1_5_1 [36] $end
$var wire 1 .5 l1_5_1 [35] $end
$var wire 1 /5 l1_5_1 [34] $end
$var wire 1 05 l1_5_1 [33] $end
$var wire 1 15 l1_5_1 [32] $end
$var wire 1 25 l1_5_1 [31] $end
$var wire 1 35 l1_5_1 [30] $end
$var wire 1 45 l1_5_1 [29] $end
$var wire 1 55 l1_5_1 [28] $end
$var wire 1 65 l1_5_1 [27] $end
$var wire 1 75 l1_5_1 [26] $end
$var wire 1 85 l1_5_1 [25] $end
$var wire 1 95 l1_5_1 [24] $end
$var wire 1 :5 l1_5_1 [23] $end
$var wire 1 ;5 l1_5_1 [22] $end
$var wire 1 <5 l1_5_1 [21] $end
$var wire 1 =5 l1_5_1 [20] $end
$var wire 1 >5 l1_5_1 [19] $end
$var wire 1 ?5 l1_5_1 [18] $end
$var wire 1 @5 l1_5_1 [17] $end
$var wire 1 A5 l1_5_1 [16] $end
$var wire 1 B5 l1_5_1 [15] $end
$var wire 1 C5 l1_5_1 [14] $end
$var wire 1 D5 l1_5_1 [13] $end
$var wire 1 E5 l1_5_1 [12] $end
$var wire 1 F5 l1_5_1 [11] $end
$var wire 1 G5 l1_5_1 [10] $end
$var wire 1 H5 l1_5_1 [9] $end
$var wire 1 I5 l1_5_1 [8] $end
$var wire 1 J5 l1_5_1 [7] $end
$var wire 1 K5 l1_5_1 [6] $end
$var wire 1 L5 l1_5_1 [5] $end
$var wire 1 M5 l1_5_1 [4] $end
$var wire 1 N5 l1_5_1 [3] $end
$var wire 1 O5 l1_5_1 [2] $end
$var wire 1 P5 l1_5_1 [1] $end
$var wire 1 Q5 l1_5_1 [0] $end
$var wire 1 R5 l1_5_2 [39] $end
$var wire 1 S5 l1_5_2 [38] $end
$var wire 1 T5 l1_5_2 [37] $end
$var wire 1 U5 l1_5_2 [36] $end
$var wire 1 V5 l1_5_2 [35] $end
$var wire 1 W5 l1_5_2 [34] $end
$var wire 1 X5 l1_5_2 [33] $end
$var wire 1 Y5 l1_5_2 [32] $end
$var wire 1 Z5 l1_5_2 [31] $end
$var wire 1 [5 l1_5_2 [30] $end
$var wire 1 \5 l1_5_2 [29] $end
$var wire 1 ]5 l1_5_2 [28] $end
$var wire 1 ^5 l1_5_2 [27] $end
$var wire 1 _5 l1_5_2 [26] $end
$var wire 1 `5 l1_5_2 [25] $end
$var wire 1 a5 l1_5_2 [24] $end
$var wire 1 b5 l1_5_2 [23] $end
$var wire 1 c5 l1_5_2 [22] $end
$var wire 1 d5 l1_5_2 [21] $end
$var wire 1 e5 l1_5_2 [20] $end
$var wire 1 f5 l1_5_2 [19] $end
$var wire 1 g5 l1_5_2 [18] $end
$var wire 1 h5 l1_5_2 [17] $end
$var wire 1 i5 l1_5_2 [16] $end
$var wire 1 j5 l1_5_2 [15] $end
$var wire 1 k5 l1_5_2 [14] $end
$var wire 1 l5 l1_5_2 [13] $end
$var wire 1 m5 l1_5_2 [12] $end
$var wire 1 n5 l1_5_2 [11] $end
$var wire 1 o5 l1_5_2 [10] $end
$var wire 1 p5 l1_5_2 [9] $end
$var wire 1 q5 l1_5_2 [8] $end
$var wire 1 r5 l1_5_2 [7] $end
$var wire 1 s5 l1_5_2 [6] $end
$var wire 1 t5 l1_5_2 [5] $end
$var wire 1 u5 l1_5_2 [4] $end
$var wire 1 v5 l1_5_2 [3] $end
$var wire 1 w5 l1_5_2 [2] $end
$var wire 1 x5 l1_5_2 [1] $end
$var wire 1 y5 l1_5_2 [0] $end
$var wire 1 z5 l1_5_cin [39] $end
$var wire 1 {5 l1_5_cin [38] $end
$var wire 1 |5 l1_5_cin [37] $end
$var wire 1 }5 l1_5_cin [36] $end
$var wire 1 ~5 l1_5_cin [35] $end
$var wire 1 !6 l1_5_cin [34] $end
$var wire 1 "6 l1_5_cin [33] $end
$var wire 1 #6 l1_5_cin [32] $end
$var wire 1 $6 l1_5_cin [31] $end
$var wire 1 %6 l1_5_cin [30] $end
$var wire 1 &6 l1_5_cin [29] $end
$var wire 1 '6 l1_5_cin [28] $end
$var wire 1 (6 l1_5_cin [27] $end
$var wire 1 )6 l1_5_cin [26] $end
$var wire 1 *6 l1_5_cin [25] $end
$var wire 1 +6 l1_5_cin [24] $end
$var wire 1 ,6 l1_5_cin [23] $end
$var wire 1 -6 l1_5_cin [22] $end
$var wire 1 .6 l1_5_cin [21] $end
$var wire 1 /6 l1_5_cin [20] $end
$var wire 1 06 l1_5_cin [19] $end
$var wire 1 16 l1_5_cin [18] $end
$var wire 1 26 l1_5_cin [17] $end
$var wire 1 36 l1_5_cin [16] $end
$var wire 1 46 l1_5_cin [15] $end
$var wire 1 56 l1_5_cin [14] $end
$var wire 1 66 l1_5_cin [13] $end
$var wire 1 76 l1_5_cin [12] $end
$var wire 1 86 l1_5_cin [11] $end
$var wire 1 96 l1_5_cin [10] $end
$var wire 1 :6 l1_5_cin [9] $end
$var wire 1 ;6 l1_5_cin [8] $end
$var wire 1 <6 l1_5_cin [7] $end
$var wire 1 =6 l1_5_cin [6] $end
$var wire 1 >6 l1_5_cin [5] $end
$var wire 1 ?6 l1_5_cin [4] $end
$var wire 1 @6 l1_5_cin [3] $end
$var wire 1 A6 l1_5_cin [2] $end
$var wire 1 B6 l1_5_cin [1] $end
$var wire 1 C6 l1_5_cin [0] $end
$var wire 1 D6 l1_5_cout [39] $end
$var wire 1 E6 l1_5_cout [38] $end
$var wire 1 F6 l1_5_cout [37] $end
$var wire 1 G6 l1_5_cout [36] $end
$var wire 1 H6 l1_5_cout [35] $end
$var wire 1 I6 l1_5_cout [34] $end
$var wire 1 J6 l1_5_cout [33] $end
$var wire 1 K6 l1_5_cout [32] $end
$var wire 1 L6 l1_5_cout [31] $end
$var wire 1 M6 l1_5_cout [30] $end
$var wire 1 N6 l1_5_cout [29] $end
$var wire 1 O6 l1_5_cout [28] $end
$var wire 1 P6 l1_5_cout [27] $end
$var wire 1 Q6 l1_5_cout [26] $end
$var wire 1 R6 l1_5_cout [25] $end
$var wire 1 S6 l1_5_cout [24] $end
$var wire 1 T6 l1_5_cout [23] $end
$var wire 1 U6 l1_5_cout [22] $end
$var wire 1 V6 l1_5_cout [21] $end
$var wire 1 W6 l1_5_cout [20] $end
$var wire 1 X6 l1_5_cout [19] $end
$var wire 1 Y6 l1_5_cout [18] $end
$var wire 1 Z6 l1_5_cout [17] $end
$var wire 1 [6 l1_5_cout [16] $end
$var wire 1 \6 l1_5_cout [15] $end
$var wire 1 ]6 l1_5_cout [14] $end
$var wire 1 ^6 l1_5_cout [13] $end
$var wire 1 _6 l1_5_cout [12] $end
$var wire 1 `6 l1_5_cout [11] $end
$var wire 1 a6 l1_5_cout [10] $end
$var wire 1 b6 l1_5_cout [9] $end
$var wire 1 c6 l1_5_cout [8] $end
$var wire 1 d6 l1_5_cout [7] $end
$var wire 1 e6 l1_5_cout [6] $end
$var wire 1 f6 l1_5_cout [5] $end
$var wire 1 g6 l1_5_cout [4] $end
$var wire 1 h6 l1_5_cout [3] $end
$var wire 1 i6 l1_5_cout [2] $end
$var wire 1 j6 l1_5_cout [1] $end
$var wire 1 k6 l1_5_cout [0] $end
$var wire 1 l6 l1_5_s [39] $end
$var wire 1 m6 l1_5_s [38] $end
$var wire 1 n6 l1_5_s [37] $end
$var wire 1 o6 l1_5_s [36] $end
$var wire 1 p6 l1_5_s [35] $end
$var wire 1 q6 l1_5_s [34] $end
$var wire 1 r6 l1_5_s [33] $end
$var wire 1 s6 l1_5_s [32] $end
$var wire 1 t6 l1_5_s [31] $end
$var wire 1 u6 l1_5_s [30] $end
$var wire 1 v6 l1_5_s [29] $end
$var wire 1 w6 l1_5_s [28] $end
$var wire 1 x6 l1_5_s [27] $end
$var wire 1 y6 l1_5_s [26] $end
$var wire 1 z6 l1_5_s [25] $end
$var wire 1 {6 l1_5_s [24] $end
$var wire 1 |6 l1_5_s [23] $end
$var wire 1 }6 l1_5_s [22] $end
$var wire 1 ~6 l1_5_s [21] $end
$var wire 1 !7 l1_5_s [20] $end
$var wire 1 "7 l1_5_s [19] $end
$var wire 1 #7 l1_5_s [18] $end
$var wire 1 $7 l1_5_s [17] $end
$var wire 1 %7 l1_5_s [16] $end
$var wire 1 &7 l1_5_s [15] $end
$var wire 1 '7 l1_5_s [14] $end
$var wire 1 (7 l1_5_s [13] $end
$var wire 1 )7 l1_5_s [12] $end
$var wire 1 *7 l1_5_s [11] $end
$var wire 1 +7 l1_5_s [10] $end
$var wire 1 ,7 l1_5_s [9] $end
$var wire 1 -7 l1_5_s [8] $end
$var wire 1 .7 l1_5_s [7] $end
$var wire 1 /7 l1_5_s [6] $end
$var wire 1 07 l1_5_s [5] $end
$var wire 1 17 l1_5_s [4] $end
$var wire 1 27 l1_5_s [3] $end
$var wire 1 37 l1_5_s [2] $end
$var wire 1 47 l1_5_s [1] $end
$var wire 1 57 l1_5_s [0] $end
$var wire 1 67 l1_5_ca [39] $end
$var wire 1 77 l1_5_ca [38] $end
$var wire 1 87 l1_5_ca [37] $end
$var wire 1 97 l1_5_ca [36] $end
$var wire 1 :7 l1_5_ca [35] $end
$var wire 1 ;7 l1_5_ca [34] $end
$var wire 1 <7 l1_5_ca [33] $end
$var wire 1 =7 l1_5_ca [32] $end
$var wire 1 >7 l1_5_ca [31] $end
$var wire 1 ?7 l1_5_ca [30] $end
$var wire 1 @7 l1_5_ca [29] $end
$var wire 1 A7 l1_5_ca [28] $end
$var wire 1 B7 l1_5_ca [27] $end
$var wire 1 C7 l1_5_ca [26] $end
$var wire 1 D7 l1_5_ca [25] $end
$var wire 1 E7 l1_5_ca [24] $end
$var wire 1 F7 l1_5_ca [23] $end
$var wire 1 G7 l1_5_ca [22] $end
$var wire 1 H7 l1_5_ca [21] $end
$var wire 1 I7 l1_5_ca [20] $end
$var wire 1 J7 l1_5_ca [19] $end
$var wire 1 K7 l1_5_ca [18] $end
$var wire 1 L7 l1_5_ca [17] $end
$var wire 1 M7 l1_5_ca [16] $end
$var wire 1 N7 l1_5_ca [15] $end
$var wire 1 O7 l1_5_ca [14] $end
$var wire 1 P7 l1_5_ca [13] $end
$var wire 1 Q7 l1_5_ca [12] $end
$var wire 1 R7 l1_5_ca [11] $end
$var wire 1 S7 l1_5_ca [10] $end
$var wire 1 T7 l1_5_ca [9] $end
$var wire 1 U7 l1_5_ca [8] $end
$var wire 1 V7 l1_5_ca [7] $end
$var wire 1 W7 l1_5_ca [6] $end
$var wire 1 X7 l1_5_ca [5] $end
$var wire 1 Y7 l1_5_ca [4] $end
$var wire 1 Z7 l1_5_ca [3] $end
$var wire 1 [7 l1_5_ca [2] $end
$var wire 1 \7 l1_5_ca [1] $end
$var wire 1 ]7 l1_5_ca [0] $end
$var wire 1 ^7 l1_6_0 [37] $end
$var wire 1 _7 l1_6_0 [36] $end
$var wire 1 `7 l1_6_0 [35] $end
$var wire 1 a7 l1_6_0 [34] $end
$var wire 1 b7 l1_6_0 [33] $end
$var wire 1 c7 l1_6_0 [32] $end
$var wire 1 d7 l1_6_0 [31] $end
$var wire 1 e7 l1_6_0 [30] $end
$var wire 1 f7 l1_6_0 [29] $end
$var wire 1 g7 l1_6_0 [28] $end
$var wire 1 h7 l1_6_0 [27] $end
$var wire 1 i7 l1_6_0 [26] $end
$var wire 1 j7 l1_6_0 [25] $end
$var wire 1 k7 l1_6_0 [24] $end
$var wire 1 l7 l1_6_0 [23] $end
$var wire 1 m7 l1_6_0 [22] $end
$var wire 1 n7 l1_6_0 [21] $end
$var wire 1 o7 l1_6_0 [20] $end
$var wire 1 p7 l1_6_0 [19] $end
$var wire 1 q7 l1_6_0 [18] $end
$var wire 1 r7 l1_6_0 [17] $end
$var wire 1 s7 l1_6_0 [16] $end
$var wire 1 t7 l1_6_0 [15] $end
$var wire 1 u7 l1_6_0 [14] $end
$var wire 1 v7 l1_6_0 [13] $end
$var wire 1 w7 l1_6_0 [12] $end
$var wire 1 x7 l1_6_0 [11] $end
$var wire 1 y7 l1_6_0 [10] $end
$var wire 1 z7 l1_6_0 [9] $end
$var wire 1 {7 l1_6_0 [8] $end
$var wire 1 |7 l1_6_0 [7] $end
$var wire 1 }7 l1_6_0 [6] $end
$var wire 1 ~7 l1_6_0 [5] $end
$var wire 1 !8 l1_6_0 [4] $end
$var wire 1 "8 l1_6_0 [3] $end
$var wire 1 #8 l1_6_0 [2] $end
$var wire 1 $8 l1_6_0 [1] $end
$var wire 1 %8 l1_6_0 [0] $end
$var wire 1 &8 l1_6_1 [37] $end
$var wire 1 '8 l1_6_1 [36] $end
$var wire 1 (8 l1_6_1 [35] $end
$var wire 1 )8 l1_6_1 [34] $end
$var wire 1 *8 l1_6_1 [33] $end
$var wire 1 +8 l1_6_1 [32] $end
$var wire 1 ,8 l1_6_1 [31] $end
$var wire 1 -8 l1_6_1 [30] $end
$var wire 1 .8 l1_6_1 [29] $end
$var wire 1 /8 l1_6_1 [28] $end
$var wire 1 08 l1_6_1 [27] $end
$var wire 1 18 l1_6_1 [26] $end
$var wire 1 28 l1_6_1 [25] $end
$var wire 1 38 l1_6_1 [24] $end
$var wire 1 48 l1_6_1 [23] $end
$var wire 1 58 l1_6_1 [22] $end
$var wire 1 68 l1_6_1 [21] $end
$var wire 1 78 l1_6_1 [20] $end
$var wire 1 88 l1_6_1 [19] $end
$var wire 1 98 l1_6_1 [18] $end
$var wire 1 :8 l1_6_1 [17] $end
$var wire 1 ;8 l1_6_1 [16] $end
$var wire 1 <8 l1_6_1 [15] $end
$var wire 1 =8 l1_6_1 [14] $end
$var wire 1 >8 l1_6_1 [13] $end
$var wire 1 ?8 l1_6_1 [12] $end
$var wire 1 @8 l1_6_1 [11] $end
$var wire 1 A8 l1_6_1 [10] $end
$var wire 1 B8 l1_6_1 [9] $end
$var wire 1 C8 l1_6_1 [8] $end
$var wire 1 D8 l1_6_1 [7] $end
$var wire 1 E8 l1_6_1 [6] $end
$var wire 1 F8 l1_6_1 [5] $end
$var wire 1 G8 l1_6_1 [4] $end
$var wire 1 H8 l1_6_1 [3] $end
$var wire 1 I8 l1_6_1 [2] $end
$var wire 1 J8 l1_6_1 [1] $end
$var wire 1 K8 l1_6_1 [0] $end
$var wire 1 L8 l1_6_2 [37] $end
$var wire 1 M8 l1_6_2 [36] $end
$var wire 1 N8 l1_6_2 [35] $end
$var wire 1 O8 l1_6_2 [34] $end
$var wire 1 P8 l1_6_2 [33] $end
$var wire 1 Q8 l1_6_2 [32] $end
$var wire 1 R8 l1_6_2 [31] $end
$var wire 1 S8 l1_6_2 [30] $end
$var wire 1 T8 l1_6_2 [29] $end
$var wire 1 U8 l1_6_2 [28] $end
$var wire 1 V8 l1_6_2 [27] $end
$var wire 1 W8 l1_6_2 [26] $end
$var wire 1 X8 l1_6_2 [25] $end
$var wire 1 Y8 l1_6_2 [24] $end
$var wire 1 Z8 l1_6_2 [23] $end
$var wire 1 [8 l1_6_2 [22] $end
$var wire 1 \8 l1_6_2 [21] $end
$var wire 1 ]8 l1_6_2 [20] $end
$var wire 1 ^8 l1_6_2 [19] $end
$var wire 1 _8 l1_6_2 [18] $end
$var wire 1 `8 l1_6_2 [17] $end
$var wire 1 a8 l1_6_2 [16] $end
$var wire 1 b8 l1_6_2 [15] $end
$var wire 1 c8 l1_6_2 [14] $end
$var wire 1 d8 l1_6_2 [13] $end
$var wire 1 e8 l1_6_2 [12] $end
$var wire 1 f8 l1_6_2 [11] $end
$var wire 1 g8 l1_6_2 [10] $end
$var wire 1 h8 l1_6_2 [9] $end
$var wire 1 i8 l1_6_2 [8] $end
$var wire 1 j8 l1_6_2 [7] $end
$var wire 1 k8 l1_6_2 [6] $end
$var wire 1 l8 l1_6_2 [5] $end
$var wire 1 m8 l1_6_2 [4] $end
$var wire 1 n8 l1_6_2 [3] $end
$var wire 1 o8 l1_6_2 [2] $end
$var wire 1 p8 l1_6_2 [1] $end
$var wire 1 q8 l1_6_2 [0] $end
$var wire 1 r8 l1_6_cin [37] $end
$var wire 1 s8 l1_6_cin [36] $end
$var wire 1 t8 l1_6_cin [35] $end
$var wire 1 u8 l1_6_cin [34] $end
$var wire 1 v8 l1_6_cin [33] $end
$var wire 1 w8 l1_6_cin [32] $end
$var wire 1 x8 l1_6_cin [31] $end
$var wire 1 y8 l1_6_cin [30] $end
$var wire 1 z8 l1_6_cin [29] $end
$var wire 1 {8 l1_6_cin [28] $end
$var wire 1 |8 l1_6_cin [27] $end
$var wire 1 }8 l1_6_cin [26] $end
$var wire 1 ~8 l1_6_cin [25] $end
$var wire 1 !9 l1_6_cin [24] $end
$var wire 1 "9 l1_6_cin [23] $end
$var wire 1 #9 l1_6_cin [22] $end
$var wire 1 $9 l1_6_cin [21] $end
$var wire 1 %9 l1_6_cin [20] $end
$var wire 1 &9 l1_6_cin [19] $end
$var wire 1 '9 l1_6_cin [18] $end
$var wire 1 (9 l1_6_cin [17] $end
$var wire 1 )9 l1_6_cin [16] $end
$var wire 1 *9 l1_6_cin [15] $end
$var wire 1 +9 l1_6_cin [14] $end
$var wire 1 ,9 l1_6_cin [13] $end
$var wire 1 -9 l1_6_cin [12] $end
$var wire 1 .9 l1_6_cin [11] $end
$var wire 1 /9 l1_6_cin [10] $end
$var wire 1 09 l1_6_cin [9] $end
$var wire 1 19 l1_6_cin [8] $end
$var wire 1 29 l1_6_cin [7] $end
$var wire 1 39 l1_6_cin [6] $end
$var wire 1 49 l1_6_cin [5] $end
$var wire 1 59 l1_6_cin [4] $end
$var wire 1 69 l1_6_cin [3] $end
$var wire 1 79 l1_6_cin [2] $end
$var wire 1 89 l1_6_cin [1] $end
$var wire 1 99 l1_6_cin [0] $end
$var wire 1 :9 l1_6_cout [37] $end
$var wire 1 ;9 l1_6_cout [36] $end
$var wire 1 <9 l1_6_cout [35] $end
$var wire 1 =9 l1_6_cout [34] $end
$var wire 1 >9 l1_6_cout [33] $end
$var wire 1 ?9 l1_6_cout [32] $end
$var wire 1 @9 l1_6_cout [31] $end
$var wire 1 A9 l1_6_cout [30] $end
$var wire 1 B9 l1_6_cout [29] $end
$var wire 1 C9 l1_6_cout [28] $end
$var wire 1 D9 l1_6_cout [27] $end
$var wire 1 E9 l1_6_cout [26] $end
$var wire 1 F9 l1_6_cout [25] $end
$var wire 1 G9 l1_6_cout [24] $end
$var wire 1 H9 l1_6_cout [23] $end
$var wire 1 I9 l1_6_cout [22] $end
$var wire 1 J9 l1_6_cout [21] $end
$var wire 1 K9 l1_6_cout [20] $end
$var wire 1 L9 l1_6_cout [19] $end
$var wire 1 M9 l1_6_cout [18] $end
$var wire 1 N9 l1_6_cout [17] $end
$var wire 1 O9 l1_6_cout [16] $end
$var wire 1 P9 l1_6_cout [15] $end
$var wire 1 Q9 l1_6_cout [14] $end
$var wire 1 R9 l1_6_cout [13] $end
$var wire 1 S9 l1_6_cout [12] $end
$var wire 1 T9 l1_6_cout [11] $end
$var wire 1 U9 l1_6_cout [10] $end
$var wire 1 V9 l1_6_cout [9] $end
$var wire 1 W9 l1_6_cout [8] $end
$var wire 1 X9 l1_6_cout [7] $end
$var wire 1 Y9 l1_6_cout [6] $end
$var wire 1 Z9 l1_6_cout [5] $end
$var wire 1 [9 l1_6_cout [4] $end
$var wire 1 \9 l1_6_cout [3] $end
$var wire 1 ]9 l1_6_cout [2] $end
$var wire 1 ^9 l1_6_cout [1] $end
$var wire 1 _9 l1_6_cout [0] $end
$var wire 1 `9 l1_6_s [37] $end
$var wire 1 a9 l1_6_s [36] $end
$var wire 1 b9 l1_6_s [35] $end
$var wire 1 c9 l1_6_s [34] $end
$var wire 1 d9 l1_6_s [33] $end
$var wire 1 e9 l1_6_s [32] $end
$var wire 1 f9 l1_6_s [31] $end
$var wire 1 g9 l1_6_s [30] $end
$var wire 1 h9 l1_6_s [29] $end
$var wire 1 i9 l1_6_s [28] $end
$var wire 1 j9 l1_6_s [27] $end
$var wire 1 k9 l1_6_s [26] $end
$var wire 1 l9 l1_6_s [25] $end
$var wire 1 m9 l1_6_s [24] $end
$var wire 1 n9 l1_6_s [23] $end
$var wire 1 o9 l1_6_s [22] $end
$var wire 1 p9 l1_6_s [21] $end
$var wire 1 q9 l1_6_s [20] $end
$var wire 1 r9 l1_6_s [19] $end
$var wire 1 s9 l1_6_s [18] $end
$var wire 1 t9 l1_6_s [17] $end
$var wire 1 u9 l1_6_s [16] $end
$var wire 1 v9 l1_6_s [15] $end
$var wire 1 w9 l1_6_s [14] $end
$var wire 1 x9 l1_6_s [13] $end
$var wire 1 y9 l1_6_s [12] $end
$var wire 1 z9 l1_6_s [11] $end
$var wire 1 {9 l1_6_s [10] $end
$var wire 1 |9 l1_6_s [9] $end
$var wire 1 }9 l1_6_s [8] $end
$var wire 1 ~9 l1_6_s [7] $end
$var wire 1 !: l1_6_s [6] $end
$var wire 1 ": l1_6_s [5] $end
$var wire 1 #: l1_6_s [4] $end
$var wire 1 $: l1_6_s [3] $end
$var wire 1 %: l1_6_s [2] $end
$var wire 1 &: l1_6_s [1] $end
$var wire 1 ': l1_6_s [0] $end
$var wire 1 (: l1_6_ca [37] $end
$var wire 1 ): l1_6_ca [36] $end
$var wire 1 *: l1_6_ca [35] $end
$var wire 1 +: l1_6_ca [34] $end
$var wire 1 ,: l1_6_ca [33] $end
$var wire 1 -: l1_6_ca [32] $end
$var wire 1 .: l1_6_ca [31] $end
$var wire 1 /: l1_6_ca [30] $end
$var wire 1 0: l1_6_ca [29] $end
$var wire 1 1: l1_6_ca [28] $end
$var wire 1 2: l1_6_ca [27] $end
$var wire 1 3: l1_6_ca [26] $end
$var wire 1 4: l1_6_ca [25] $end
$var wire 1 5: l1_6_ca [24] $end
$var wire 1 6: l1_6_ca [23] $end
$var wire 1 7: l1_6_ca [22] $end
$var wire 1 8: l1_6_ca [21] $end
$var wire 1 9: l1_6_ca [20] $end
$var wire 1 :: l1_6_ca [19] $end
$var wire 1 ;: l1_6_ca [18] $end
$var wire 1 <: l1_6_ca [17] $end
$var wire 1 =: l1_6_ca [16] $end
$var wire 1 >: l1_6_ca [15] $end
$var wire 1 ?: l1_6_ca [14] $end
$var wire 1 @: l1_6_ca [13] $end
$var wire 1 A: l1_6_ca [12] $end
$var wire 1 B: l1_6_ca [11] $end
$var wire 1 C: l1_6_ca [10] $end
$var wire 1 D: l1_6_ca [9] $end
$var wire 1 E: l1_6_ca [8] $end
$var wire 1 F: l1_6_ca [7] $end
$var wire 1 G: l1_6_ca [6] $end
$var wire 1 H: l1_6_ca [5] $end
$var wire 1 I: l1_6_ca [4] $end
$var wire 1 J: l1_6_ca [3] $end
$var wire 1 K: l1_6_ca [2] $end
$var wire 1 L: l1_6_ca [1] $end
$var wire 1 M: l1_6_ca [0] $end
$var reg 36 N: l1_s1_reg [35:0] $end
$var reg 36 O: l1_c1_reg [35:0] $end
$var reg 40 P: l1_s2_reg [39:0] $end
$var reg 40 Q: l1_c2_reg [39:0] $end
$var reg 40 R: l1_s3_reg [39:0] $end
$var reg 40 S: l1_c3_reg [39:0] $end
$var reg 40 T: l1_s4_reg [39:0] $end
$var reg 40 U: l1_c4_reg [39:0] $end
$var reg 40 V: l1_s5_reg [39:0] $end
$var reg 40 W: l1_c5_reg [39:0] $end
$var reg 38 X: l1_s6_reg [37:0] $end
$var reg 38 Y: l1_c6_reg [37:0] $end
$var wire 1 Z: l2_1_0 [42] $end
$var wire 1 [: l2_1_0 [41] $end
$var wire 1 \: l2_1_0 [40] $end
$var wire 1 ]: l2_1_0 [39] $end
$var wire 1 ^: l2_1_0 [38] $end
$var wire 1 _: l2_1_0 [37] $end
$var wire 1 `: l2_1_0 [36] $end
$var wire 1 a: l2_1_0 [35] $end
$var wire 1 b: l2_1_0 [34] $end
$var wire 1 c: l2_1_0 [33] $end
$var wire 1 d: l2_1_0 [32] $end
$var wire 1 e: l2_1_0 [31] $end
$var wire 1 f: l2_1_0 [30] $end
$var wire 1 g: l2_1_0 [29] $end
$var wire 1 h: l2_1_0 [28] $end
$var wire 1 i: l2_1_0 [27] $end
$var wire 1 j: l2_1_0 [26] $end
$var wire 1 k: l2_1_0 [25] $end
$var wire 1 l: l2_1_0 [24] $end
$var wire 1 m: l2_1_0 [23] $end
$var wire 1 n: l2_1_0 [22] $end
$var wire 1 o: l2_1_0 [21] $end
$var wire 1 p: l2_1_0 [20] $end
$var wire 1 q: l2_1_0 [19] $end
$var wire 1 r: l2_1_0 [18] $end
$var wire 1 s: l2_1_0 [17] $end
$var wire 1 t: l2_1_0 [16] $end
$var wire 1 u: l2_1_0 [15] $end
$var wire 1 v: l2_1_0 [14] $end
$var wire 1 w: l2_1_0 [13] $end
$var wire 1 x: l2_1_0 [12] $end
$var wire 1 y: l2_1_0 [11] $end
$var wire 1 z: l2_1_0 [10] $end
$var wire 1 {: l2_1_0 [9] $end
$var wire 1 |: l2_1_0 [8] $end
$var wire 1 }: l2_1_0 [7] $end
$var wire 1 ~: l2_1_0 [6] $end
$var wire 1 !; l2_1_0 [5] $end
$var wire 1 "; l2_1_0 [4] $end
$var wire 1 #; l2_1_0 [3] $end
$var wire 1 $; l2_1_0 [2] $end
$var wire 1 %; l2_1_0 [1] $end
$var wire 1 &; l2_1_0 [0] $end
$var wire 1 '; l2_1_1 [42] $end
$var wire 1 (; l2_1_1 [41] $end
$var wire 1 ); l2_1_1 [40] $end
$var wire 1 *; l2_1_1 [39] $end
$var wire 1 +; l2_1_1 [38] $end
$var wire 1 ,; l2_1_1 [37] $end
$var wire 1 -; l2_1_1 [36] $end
$var wire 1 .; l2_1_1 [35] $end
$var wire 1 /; l2_1_1 [34] $end
$var wire 1 0; l2_1_1 [33] $end
$var wire 1 1; l2_1_1 [32] $end
$var wire 1 2; l2_1_1 [31] $end
$var wire 1 3; l2_1_1 [30] $end
$var wire 1 4; l2_1_1 [29] $end
$var wire 1 5; l2_1_1 [28] $end
$var wire 1 6; l2_1_1 [27] $end
$var wire 1 7; l2_1_1 [26] $end
$var wire 1 8; l2_1_1 [25] $end
$var wire 1 9; l2_1_1 [24] $end
$var wire 1 :; l2_1_1 [23] $end
$var wire 1 ;; l2_1_1 [22] $end
$var wire 1 <; l2_1_1 [21] $end
$var wire 1 =; l2_1_1 [20] $end
$var wire 1 >; l2_1_1 [19] $end
$var wire 1 ?; l2_1_1 [18] $end
$var wire 1 @; l2_1_1 [17] $end
$var wire 1 A; l2_1_1 [16] $end
$var wire 1 B; l2_1_1 [15] $end
$var wire 1 C; l2_1_1 [14] $end
$var wire 1 D; l2_1_1 [13] $end
$var wire 1 E; l2_1_1 [12] $end
$var wire 1 F; l2_1_1 [11] $end
$var wire 1 G; l2_1_1 [10] $end
$var wire 1 H; l2_1_1 [9] $end
$var wire 1 I; l2_1_1 [8] $end
$var wire 1 J; l2_1_1 [7] $end
$var wire 1 K; l2_1_1 [6] $end
$var wire 1 L; l2_1_1 [5] $end
$var wire 1 M; l2_1_1 [4] $end
$var wire 1 N; l2_1_1 [3] $end
$var wire 1 O; l2_1_1 [2] $end
$var wire 1 P; l2_1_1 [1] $end
$var wire 1 Q; l2_1_1 [0] $end
$var wire 1 R; l2_1_2 [42] $end
$var wire 1 S; l2_1_2 [41] $end
$var wire 1 T; l2_1_2 [40] $end
$var wire 1 U; l2_1_2 [39] $end
$var wire 1 V; l2_1_2 [38] $end
$var wire 1 W; l2_1_2 [37] $end
$var wire 1 X; l2_1_2 [36] $end
$var wire 1 Y; l2_1_2 [35] $end
$var wire 1 Z; l2_1_2 [34] $end
$var wire 1 [; l2_1_2 [33] $end
$var wire 1 \; l2_1_2 [32] $end
$var wire 1 ]; l2_1_2 [31] $end
$var wire 1 ^; l2_1_2 [30] $end
$var wire 1 _; l2_1_2 [29] $end
$var wire 1 `; l2_1_2 [28] $end
$var wire 1 a; l2_1_2 [27] $end
$var wire 1 b; l2_1_2 [26] $end
$var wire 1 c; l2_1_2 [25] $end
$var wire 1 d; l2_1_2 [24] $end
$var wire 1 e; l2_1_2 [23] $end
$var wire 1 f; l2_1_2 [22] $end
$var wire 1 g; l2_1_2 [21] $end
$var wire 1 h; l2_1_2 [20] $end
$var wire 1 i; l2_1_2 [19] $end
$var wire 1 j; l2_1_2 [18] $end
$var wire 1 k; l2_1_2 [17] $end
$var wire 1 l; l2_1_2 [16] $end
$var wire 1 m; l2_1_2 [15] $end
$var wire 1 n; l2_1_2 [14] $end
$var wire 1 o; l2_1_2 [13] $end
$var wire 1 p; l2_1_2 [12] $end
$var wire 1 q; l2_1_2 [11] $end
$var wire 1 r; l2_1_2 [10] $end
$var wire 1 s; l2_1_2 [9] $end
$var wire 1 t; l2_1_2 [8] $end
$var wire 1 u; l2_1_2 [7] $end
$var wire 1 v; l2_1_2 [6] $end
$var wire 1 w; l2_1_2 [5] $end
$var wire 1 x; l2_1_2 [4] $end
$var wire 1 y; l2_1_2 [3] $end
$var wire 1 z; l2_1_2 [2] $end
$var wire 1 {; l2_1_2 [1] $end
$var wire 1 |; l2_1_2 [0] $end
$var wire 1 }; l2_1_3 [42] $end
$var wire 1 ~; l2_1_3 [41] $end
$var wire 1 !< l2_1_3 [40] $end
$var wire 1 "< l2_1_3 [39] $end
$var wire 1 #< l2_1_3 [38] $end
$var wire 1 $< l2_1_3 [37] $end
$var wire 1 %< l2_1_3 [36] $end
$var wire 1 &< l2_1_3 [35] $end
$var wire 1 '< l2_1_3 [34] $end
$var wire 1 (< l2_1_3 [33] $end
$var wire 1 )< l2_1_3 [32] $end
$var wire 1 *< l2_1_3 [31] $end
$var wire 1 +< l2_1_3 [30] $end
$var wire 1 ,< l2_1_3 [29] $end
$var wire 1 -< l2_1_3 [28] $end
$var wire 1 .< l2_1_3 [27] $end
$var wire 1 /< l2_1_3 [26] $end
$var wire 1 0< l2_1_3 [25] $end
$var wire 1 1< l2_1_3 [24] $end
$var wire 1 2< l2_1_3 [23] $end
$var wire 1 3< l2_1_3 [22] $end
$var wire 1 4< l2_1_3 [21] $end
$var wire 1 5< l2_1_3 [20] $end
$var wire 1 6< l2_1_3 [19] $end
$var wire 1 7< l2_1_3 [18] $end
$var wire 1 8< l2_1_3 [17] $end
$var wire 1 9< l2_1_3 [16] $end
$var wire 1 :< l2_1_3 [15] $end
$var wire 1 ;< l2_1_3 [14] $end
$var wire 1 << l2_1_3 [13] $end
$var wire 1 =< l2_1_3 [12] $end
$var wire 1 >< l2_1_3 [11] $end
$var wire 1 ?< l2_1_3 [10] $end
$var wire 1 @< l2_1_3 [9] $end
$var wire 1 A< l2_1_3 [8] $end
$var wire 1 B< l2_1_3 [7] $end
$var wire 1 C< l2_1_3 [6] $end
$var wire 1 D< l2_1_3 [5] $end
$var wire 1 E< l2_1_3 [4] $end
$var wire 1 F< l2_1_3 [3] $end
$var wire 1 G< l2_1_3 [2] $end
$var wire 1 H< l2_1_3 [1] $end
$var wire 1 I< l2_1_3 [0] $end
$var wire 1 J< l2_1_cin [42] $end
$var wire 1 K< l2_1_cin [41] $end
$var wire 1 L< l2_1_cin [40] $end
$var wire 1 M< l2_1_cin [39] $end
$var wire 1 N< l2_1_cin [38] $end
$var wire 1 O< l2_1_cin [37] $end
$var wire 1 P< l2_1_cin [36] $end
$var wire 1 Q< l2_1_cin [35] $end
$var wire 1 R< l2_1_cin [34] $end
$var wire 1 S< l2_1_cin [33] $end
$var wire 1 T< l2_1_cin [32] $end
$var wire 1 U< l2_1_cin [31] $end
$var wire 1 V< l2_1_cin [30] $end
$var wire 1 W< l2_1_cin [29] $end
$var wire 1 X< l2_1_cin [28] $end
$var wire 1 Y< l2_1_cin [27] $end
$var wire 1 Z< l2_1_cin [26] $end
$var wire 1 [< l2_1_cin [25] $end
$var wire 1 \< l2_1_cin [24] $end
$var wire 1 ]< l2_1_cin [23] $end
$var wire 1 ^< l2_1_cin [22] $end
$var wire 1 _< l2_1_cin [21] $end
$var wire 1 `< l2_1_cin [20] $end
$var wire 1 a< l2_1_cin [19] $end
$var wire 1 b< l2_1_cin [18] $end
$var wire 1 c< l2_1_cin [17] $end
$var wire 1 d< l2_1_cin [16] $end
$var wire 1 e< l2_1_cin [15] $end
$var wire 1 f< l2_1_cin [14] $end
$var wire 1 g< l2_1_cin [13] $end
$var wire 1 h< l2_1_cin [12] $end
$var wire 1 i< l2_1_cin [11] $end
$var wire 1 j< l2_1_cin [10] $end
$var wire 1 k< l2_1_cin [9] $end
$var wire 1 l< l2_1_cin [8] $end
$var wire 1 m< l2_1_cin [7] $end
$var wire 1 n< l2_1_cin [6] $end
$var wire 1 o< l2_1_cin [5] $end
$var wire 1 p< l2_1_cin [4] $end
$var wire 1 q< l2_1_cin [3] $end
$var wire 1 r< l2_1_cin [2] $end
$var wire 1 s< l2_1_cin [1] $end
$var wire 1 t< l2_1_cin [0] $end
$var wire 1 u< l2_1_cout [42] $end
$var wire 1 v< l2_1_cout [41] $end
$var wire 1 w< l2_1_cout [40] $end
$var wire 1 x< l2_1_cout [39] $end
$var wire 1 y< l2_1_cout [38] $end
$var wire 1 z< l2_1_cout [37] $end
$var wire 1 {< l2_1_cout [36] $end
$var wire 1 |< l2_1_cout [35] $end
$var wire 1 }< l2_1_cout [34] $end
$var wire 1 ~< l2_1_cout [33] $end
$var wire 1 != l2_1_cout [32] $end
$var wire 1 "= l2_1_cout [31] $end
$var wire 1 #= l2_1_cout [30] $end
$var wire 1 $= l2_1_cout [29] $end
$var wire 1 %= l2_1_cout [28] $end
$var wire 1 &= l2_1_cout [27] $end
$var wire 1 '= l2_1_cout [26] $end
$var wire 1 (= l2_1_cout [25] $end
$var wire 1 )= l2_1_cout [24] $end
$var wire 1 *= l2_1_cout [23] $end
$var wire 1 += l2_1_cout [22] $end
$var wire 1 ,= l2_1_cout [21] $end
$var wire 1 -= l2_1_cout [20] $end
$var wire 1 .= l2_1_cout [19] $end
$var wire 1 /= l2_1_cout [18] $end
$var wire 1 0= l2_1_cout [17] $end
$var wire 1 1= l2_1_cout [16] $end
$var wire 1 2= l2_1_cout [15] $end
$var wire 1 3= l2_1_cout [14] $end
$var wire 1 4= l2_1_cout [13] $end
$var wire 1 5= l2_1_cout [12] $end
$var wire 1 6= l2_1_cout [11] $end
$var wire 1 7= l2_1_cout [10] $end
$var wire 1 8= l2_1_cout [9] $end
$var wire 1 9= l2_1_cout [8] $end
$var wire 1 := l2_1_cout [7] $end
$var wire 1 ;= l2_1_cout [6] $end
$var wire 1 <= l2_1_cout [5] $end
$var wire 1 == l2_1_cout [4] $end
$var wire 1 >= l2_1_cout [3] $end
$var wire 1 ?= l2_1_cout [2] $end
$var wire 1 @= l2_1_cout [1] $end
$var wire 1 A= l2_1_cout [0] $end
$var wire 1 B= l2_1_s [42] $end
$var wire 1 C= l2_1_s [41] $end
$var wire 1 D= l2_1_s [40] $end
$var wire 1 E= l2_1_s [39] $end
$var wire 1 F= l2_1_s [38] $end
$var wire 1 G= l2_1_s [37] $end
$var wire 1 H= l2_1_s [36] $end
$var wire 1 I= l2_1_s [35] $end
$var wire 1 J= l2_1_s [34] $end
$var wire 1 K= l2_1_s [33] $end
$var wire 1 L= l2_1_s [32] $end
$var wire 1 M= l2_1_s [31] $end
$var wire 1 N= l2_1_s [30] $end
$var wire 1 O= l2_1_s [29] $end
$var wire 1 P= l2_1_s [28] $end
$var wire 1 Q= l2_1_s [27] $end
$var wire 1 R= l2_1_s [26] $end
$var wire 1 S= l2_1_s [25] $end
$var wire 1 T= l2_1_s [24] $end
$var wire 1 U= l2_1_s [23] $end
$var wire 1 V= l2_1_s [22] $end
$var wire 1 W= l2_1_s [21] $end
$var wire 1 X= l2_1_s [20] $end
$var wire 1 Y= l2_1_s [19] $end
$var wire 1 Z= l2_1_s [18] $end
$var wire 1 [= l2_1_s [17] $end
$var wire 1 \= l2_1_s [16] $end
$var wire 1 ]= l2_1_s [15] $end
$var wire 1 ^= l2_1_s [14] $end
$var wire 1 _= l2_1_s [13] $end
$var wire 1 `= l2_1_s [12] $end
$var wire 1 a= l2_1_s [11] $end
$var wire 1 b= l2_1_s [10] $end
$var wire 1 c= l2_1_s [9] $end
$var wire 1 d= l2_1_s [8] $end
$var wire 1 e= l2_1_s [7] $end
$var wire 1 f= l2_1_s [6] $end
$var wire 1 g= l2_1_s [5] $end
$var wire 1 h= l2_1_s [4] $end
$var wire 1 i= l2_1_s [3] $end
$var wire 1 j= l2_1_s [2] $end
$var wire 1 k= l2_1_s [1] $end
$var wire 1 l= l2_1_s [0] $end
$var wire 1 m= l2_1_ca [42] $end
$var wire 1 n= l2_1_ca [41] $end
$var wire 1 o= l2_1_ca [40] $end
$var wire 1 p= l2_1_ca [39] $end
$var wire 1 q= l2_1_ca [38] $end
$var wire 1 r= l2_1_ca [37] $end
$var wire 1 s= l2_1_ca [36] $end
$var wire 1 t= l2_1_ca [35] $end
$var wire 1 u= l2_1_ca [34] $end
$var wire 1 v= l2_1_ca [33] $end
$var wire 1 w= l2_1_ca [32] $end
$var wire 1 x= l2_1_ca [31] $end
$var wire 1 y= l2_1_ca [30] $end
$var wire 1 z= l2_1_ca [29] $end
$var wire 1 {= l2_1_ca [28] $end
$var wire 1 |= l2_1_ca [27] $end
$var wire 1 }= l2_1_ca [26] $end
$var wire 1 ~= l2_1_ca [25] $end
$var wire 1 !> l2_1_ca [24] $end
$var wire 1 "> l2_1_ca [23] $end
$var wire 1 #> l2_1_ca [22] $end
$var wire 1 $> l2_1_ca [21] $end
$var wire 1 %> l2_1_ca [20] $end
$var wire 1 &> l2_1_ca [19] $end
$var wire 1 '> l2_1_ca [18] $end
$var wire 1 (> l2_1_ca [17] $end
$var wire 1 )> l2_1_ca [16] $end
$var wire 1 *> l2_1_ca [15] $end
$var wire 1 +> l2_1_ca [14] $end
$var wire 1 ,> l2_1_ca [13] $end
$var wire 1 -> l2_1_ca [12] $end
$var wire 1 .> l2_1_ca [11] $end
$var wire 1 /> l2_1_ca [10] $end
$var wire 1 0> l2_1_ca [9] $end
$var wire 1 1> l2_1_ca [8] $end
$var wire 1 2> l2_1_ca [7] $end
$var wire 1 3> l2_1_ca [6] $end
$var wire 1 4> l2_1_ca [5] $end
$var wire 1 5> l2_1_ca [4] $end
$var wire 1 6> l2_1_ca [3] $end
$var wire 1 7> l2_1_ca [2] $end
$var wire 1 8> l2_1_ca [1] $end
$var wire 1 9> l2_1_ca [0] $end
$var wire 1 :> l2_2_0 [46] $end
$var wire 1 ;> l2_2_0 [45] $end
$var wire 1 <> l2_2_0 [44] $end
$var wire 1 => l2_2_0 [43] $end
$var wire 1 >> l2_2_0 [42] $end
$var wire 1 ?> l2_2_0 [41] $end
$var wire 1 @> l2_2_0 [40] $end
$var wire 1 A> l2_2_0 [39] $end
$var wire 1 B> l2_2_0 [38] $end
$var wire 1 C> l2_2_0 [37] $end
$var wire 1 D> l2_2_0 [36] $end
$var wire 1 E> l2_2_0 [35] $end
$var wire 1 F> l2_2_0 [34] $end
$var wire 1 G> l2_2_0 [33] $end
$var wire 1 H> l2_2_0 [32] $end
$var wire 1 I> l2_2_0 [31] $end
$var wire 1 J> l2_2_0 [30] $end
$var wire 1 K> l2_2_0 [29] $end
$var wire 1 L> l2_2_0 [28] $end
$var wire 1 M> l2_2_0 [27] $end
$var wire 1 N> l2_2_0 [26] $end
$var wire 1 O> l2_2_0 [25] $end
$var wire 1 P> l2_2_0 [24] $end
$var wire 1 Q> l2_2_0 [23] $end
$var wire 1 R> l2_2_0 [22] $end
$var wire 1 S> l2_2_0 [21] $end
$var wire 1 T> l2_2_0 [20] $end
$var wire 1 U> l2_2_0 [19] $end
$var wire 1 V> l2_2_0 [18] $end
$var wire 1 W> l2_2_0 [17] $end
$var wire 1 X> l2_2_0 [16] $end
$var wire 1 Y> l2_2_0 [15] $end
$var wire 1 Z> l2_2_0 [14] $end
$var wire 1 [> l2_2_0 [13] $end
$var wire 1 \> l2_2_0 [12] $end
$var wire 1 ]> l2_2_0 [11] $end
$var wire 1 ^> l2_2_0 [10] $end
$var wire 1 _> l2_2_0 [9] $end
$var wire 1 `> l2_2_0 [8] $end
$var wire 1 a> l2_2_0 [7] $end
$var wire 1 b> l2_2_0 [6] $end
$var wire 1 c> l2_2_0 [5] $end
$var wire 1 d> l2_2_0 [4] $end
$var wire 1 e> l2_2_0 [3] $end
$var wire 1 f> l2_2_0 [2] $end
$var wire 1 g> l2_2_0 [1] $end
$var wire 1 h> l2_2_0 [0] $end
$var wire 1 i> l2_2_1 [46] $end
$var wire 1 j> l2_2_1 [45] $end
$var wire 1 k> l2_2_1 [44] $end
$var wire 1 l> l2_2_1 [43] $end
$var wire 1 m> l2_2_1 [42] $end
$var wire 1 n> l2_2_1 [41] $end
$var wire 1 o> l2_2_1 [40] $end
$var wire 1 p> l2_2_1 [39] $end
$var wire 1 q> l2_2_1 [38] $end
$var wire 1 r> l2_2_1 [37] $end
$var wire 1 s> l2_2_1 [36] $end
$var wire 1 t> l2_2_1 [35] $end
$var wire 1 u> l2_2_1 [34] $end
$var wire 1 v> l2_2_1 [33] $end
$var wire 1 w> l2_2_1 [32] $end
$var wire 1 x> l2_2_1 [31] $end
$var wire 1 y> l2_2_1 [30] $end
$var wire 1 z> l2_2_1 [29] $end
$var wire 1 {> l2_2_1 [28] $end
$var wire 1 |> l2_2_1 [27] $end
$var wire 1 }> l2_2_1 [26] $end
$var wire 1 ~> l2_2_1 [25] $end
$var wire 1 !? l2_2_1 [24] $end
$var wire 1 "? l2_2_1 [23] $end
$var wire 1 #? l2_2_1 [22] $end
$var wire 1 $? l2_2_1 [21] $end
$var wire 1 %? l2_2_1 [20] $end
$var wire 1 &? l2_2_1 [19] $end
$var wire 1 '? l2_2_1 [18] $end
$var wire 1 (? l2_2_1 [17] $end
$var wire 1 )? l2_2_1 [16] $end
$var wire 1 *? l2_2_1 [15] $end
$var wire 1 +? l2_2_1 [14] $end
$var wire 1 ,? l2_2_1 [13] $end
$var wire 1 -? l2_2_1 [12] $end
$var wire 1 .? l2_2_1 [11] $end
$var wire 1 /? l2_2_1 [10] $end
$var wire 1 0? l2_2_1 [9] $end
$var wire 1 1? l2_2_1 [8] $end
$var wire 1 2? l2_2_1 [7] $end
$var wire 1 3? l2_2_1 [6] $end
$var wire 1 4? l2_2_1 [5] $end
$var wire 1 5? l2_2_1 [4] $end
$var wire 1 6? l2_2_1 [3] $end
$var wire 1 7? l2_2_1 [2] $end
$var wire 1 8? l2_2_1 [1] $end
$var wire 1 9? l2_2_1 [0] $end
$var wire 1 :? l2_2_2 [46] $end
$var wire 1 ;? l2_2_2 [45] $end
$var wire 1 <? l2_2_2 [44] $end
$var wire 1 =? l2_2_2 [43] $end
$var wire 1 >? l2_2_2 [42] $end
$var wire 1 ?? l2_2_2 [41] $end
$var wire 1 @? l2_2_2 [40] $end
$var wire 1 A? l2_2_2 [39] $end
$var wire 1 B? l2_2_2 [38] $end
$var wire 1 C? l2_2_2 [37] $end
$var wire 1 D? l2_2_2 [36] $end
$var wire 1 E? l2_2_2 [35] $end
$var wire 1 F? l2_2_2 [34] $end
$var wire 1 G? l2_2_2 [33] $end
$var wire 1 H? l2_2_2 [32] $end
$var wire 1 I? l2_2_2 [31] $end
$var wire 1 J? l2_2_2 [30] $end
$var wire 1 K? l2_2_2 [29] $end
$var wire 1 L? l2_2_2 [28] $end
$var wire 1 M? l2_2_2 [27] $end
$var wire 1 N? l2_2_2 [26] $end
$var wire 1 O? l2_2_2 [25] $end
$var wire 1 P? l2_2_2 [24] $end
$var wire 1 Q? l2_2_2 [23] $end
$var wire 1 R? l2_2_2 [22] $end
$var wire 1 S? l2_2_2 [21] $end
$var wire 1 T? l2_2_2 [20] $end
$var wire 1 U? l2_2_2 [19] $end
$var wire 1 V? l2_2_2 [18] $end
$var wire 1 W? l2_2_2 [17] $end
$var wire 1 X? l2_2_2 [16] $end
$var wire 1 Y? l2_2_2 [15] $end
$var wire 1 Z? l2_2_2 [14] $end
$var wire 1 [? l2_2_2 [13] $end
$var wire 1 \? l2_2_2 [12] $end
$var wire 1 ]? l2_2_2 [11] $end
$var wire 1 ^? l2_2_2 [10] $end
$var wire 1 _? l2_2_2 [9] $end
$var wire 1 `? l2_2_2 [8] $end
$var wire 1 a? l2_2_2 [7] $end
$var wire 1 b? l2_2_2 [6] $end
$var wire 1 c? l2_2_2 [5] $end
$var wire 1 d? l2_2_2 [4] $end
$var wire 1 e? l2_2_2 [3] $end
$var wire 1 f? l2_2_2 [2] $end
$var wire 1 g? l2_2_2 [1] $end
$var wire 1 h? l2_2_2 [0] $end
$var wire 1 i? l2_2_3 [46] $end
$var wire 1 j? l2_2_3 [45] $end
$var wire 1 k? l2_2_3 [44] $end
$var wire 1 l? l2_2_3 [43] $end
$var wire 1 m? l2_2_3 [42] $end
$var wire 1 n? l2_2_3 [41] $end
$var wire 1 o? l2_2_3 [40] $end
$var wire 1 p? l2_2_3 [39] $end
$var wire 1 q? l2_2_3 [38] $end
$var wire 1 r? l2_2_3 [37] $end
$var wire 1 s? l2_2_3 [36] $end
$var wire 1 t? l2_2_3 [35] $end
$var wire 1 u? l2_2_3 [34] $end
$var wire 1 v? l2_2_3 [33] $end
$var wire 1 w? l2_2_3 [32] $end
$var wire 1 x? l2_2_3 [31] $end
$var wire 1 y? l2_2_3 [30] $end
$var wire 1 z? l2_2_3 [29] $end
$var wire 1 {? l2_2_3 [28] $end
$var wire 1 |? l2_2_3 [27] $end
$var wire 1 }? l2_2_3 [26] $end
$var wire 1 ~? l2_2_3 [25] $end
$var wire 1 !@ l2_2_3 [24] $end
$var wire 1 "@ l2_2_3 [23] $end
$var wire 1 #@ l2_2_3 [22] $end
$var wire 1 $@ l2_2_3 [21] $end
$var wire 1 %@ l2_2_3 [20] $end
$var wire 1 &@ l2_2_3 [19] $end
$var wire 1 '@ l2_2_3 [18] $end
$var wire 1 (@ l2_2_3 [17] $end
$var wire 1 )@ l2_2_3 [16] $end
$var wire 1 *@ l2_2_3 [15] $end
$var wire 1 +@ l2_2_3 [14] $end
$var wire 1 ,@ l2_2_3 [13] $end
$var wire 1 -@ l2_2_3 [12] $end
$var wire 1 .@ l2_2_3 [11] $end
$var wire 1 /@ l2_2_3 [10] $end
$var wire 1 0@ l2_2_3 [9] $end
$var wire 1 1@ l2_2_3 [8] $end
$var wire 1 2@ l2_2_3 [7] $end
$var wire 1 3@ l2_2_3 [6] $end
$var wire 1 4@ l2_2_3 [5] $end
$var wire 1 5@ l2_2_3 [4] $end
$var wire 1 6@ l2_2_3 [3] $end
$var wire 1 7@ l2_2_3 [2] $end
$var wire 1 8@ l2_2_3 [1] $end
$var wire 1 9@ l2_2_3 [0] $end
$var wire 1 :@ l2_2_cin [46] $end
$var wire 1 ;@ l2_2_cin [45] $end
$var wire 1 <@ l2_2_cin [44] $end
$var wire 1 =@ l2_2_cin [43] $end
$var wire 1 >@ l2_2_cin [42] $end
$var wire 1 ?@ l2_2_cin [41] $end
$var wire 1 @@ l2_2_cin [40] $end
$var wire 1 A@ l2_2_cin [39] $end
$var wire 1 B@ l2_2_cin [38] $end
$var wire 1 C@ l2_2_cin [37] $end
$var wire 1 D@ l2_2_cin [36] $end
$var wire 1 E@ l2_2_cin [35] $end
$var wire 1 F@ l2_2_cin [34] $end
$var wire 1 G@ l2_2_cin [33] $end
$var wire 1 H@ l2_2_cin [32] $end
$var wire 1 I@ l2_2_cin [31] $end
$var wire 1 J@ l2_2_cin [30] $end
$var wire 1 K@ l2_2_cin [29] $end
$var wire 1 L@ l2_2_cin [28] $end
$var wire 1 M@ l2_2_cin [27] $end
$var wire 1 N@ l2_2_cin [26] $end
$var wire 1 O@ l2_2_cin [25] $end
$var wire 1 P@ l2_2_cin [24] $end
$var wire 1 Q@ l2_2_cin [23] $end
$var wire 1 R@ l2_2_cin [22] $end
$var wire 1 S@ l2_2_cin [21] $end
$var wire 1 T@ l2_2_cin [20] $end
$var wire 1 U@ l2_2_cin [19] $end
$var wire 1 V@ l2_2_cin [18] $end
$var wire 1 W@ l2_2_cin [17] $end
$var wire 1 X@ l2_2_cin [16] $end
$var wire 1 Y@ l2_2_cin [15] $end
$var wire 1 Z@ l2_2_cin [14] $end
$var wire 1 [@ l2_2_cin [13] $end
$var wire 1 \@ l2_2_cin [12] $end
$var wire 1 ]@ l2_2_cin [11] $end
$var wire 1 ^@ l2_2_cin [10] $end
$var wire 1 _@ l2_2_cin [9] $end
$var wire 1 `@ l2_2_cin [8] $end
$var wire 1 a@ l2_2_cin [7] $end
$var wire 1 b@ l2_2_cin [6] $end
$var wire 1 c@ l2_2_cin [5] $end
$var wire 1 d@ l2_2_cin [4] $end
$var wire 1 e@ l2_2_cin [3] $end
$var wire 1 f@ l2_2_cin [2] $end
$var wire 1 g@ l2_2_cin [1] $end
$var wire 1 h@ l2_2_cin [0] $end
$var wire 1 i@ l2_2_cout [46] $end
$var wire 1 j@ l2_2_cout [45] $end
$var wire 1 k@ l2_2_cout [44] $end
$var wire 1 l@ l2_2_cout [43] $end
$var wire 1 m@ l2_2_cout [42] $end
$var wire 1 n@ l2_2_cout [41] $end
$var wire 1 o@ l2_2_cout [40] $end
$var wire 1 p@ l2_2_cout [39] $end
$var wire 1 q@ l2_2_cout [38] $end
$var wire 1 r@ l2_2_cout [37] $end
$var wire 1 s@ l2_2_cout [36] $end
$var wire 1 t@ l2_2_cout [35] $end
$var wire 1 u@ l2_2_cout [34] $end
$var wire 1 v@ l2_2_cout [33] $end
$var wire 1 w@ l2_2_cout [32] $end
$var wire 1 x@ l2_2_cout [31] $end
$var wire 1 y@ l2_2_cout [30] $end
$var wire 1 z@ l2_2_cout [29] $end
$var wire 1 {@ l2_2_cout [28] $end
$var wire 1 |@ l2_2_cout [27] $end
$var wire 1 }@ l2_2_cout [26] $end
$var wire 1 ~@ l2_2_cout [25] $end
$var wire 1 !A l2_2_cout [24] $end
$var wire 1 "A l2_2_cout [23] $end
$var wire 1 #A l2_2_cout [22] $end
$var wire 1 $A l2_2_cout [21] $end
$var wire 1 %A l2_2_cout [20] $end
$var wire 1 &A l2_2_cout [19] $end
$var wire 1 'A l2_2_cout [18] $end
$var wire 1 (A l2_2_cout [17] $end
$var wire 1 )A l2_2_cout [16] $end
$var wire 1 *A l2_2_cout [15] $end
$var wire 1 +A l2_2_cout [14] $end
$var wire 1 ,A l2_2_cout [13] $end
$var wire 1 -A l2_2_cout [12] $end
$var wire 1 .A l2_2_cout [11] $end
$var wire 1 /A l2_2_cout [10] $end
$var wire 1 0A l2_2_cout [9] $end
$var wire 1 1A l2_2_cout [8] $end
$var wire 1 2A l2_2_cout [7] $end
$var wire 1 3A l2_2_cout [6] $end
$var wire 1 4A l2_2_cout [5] $end
$var wire 1 5A l2_2_cout [4] $end
$var wire 1 6A l2_2_cout [3] $end
$var wire 1 7A l2_2_cout [2] $end
$var wire 1 8A l2_2_cout [1] $end
$var wire 1 9A l2_2_cout [0] $end
$var wire 1 :A l2_2_s [46] $end
$var wire 1 ;A l2_2_s [45] $end
$var wire 1 <A l2_2_s [44] $end
$var wire 1 =A l2_2_s [43] $end
$var wire 1 >A l2_2_s [42] $end
$var wire 1 ?A l2_2_s [41] $end
$var wire 1 @A l2_2_s [40] $end
$var wire 1 AA l2_2_s [39] $end
$var wire 1 BA l2_2_s [38] $end
$var wire 1 CA l2_2_s [37] $end
$var wire 1 DA l2_2_s [36] $end
$var wire 1 EA l2_2_s [35] $end
$var wire 1 FA l2_2_s [34] $end
$var wire 1 GA l2_2_s [33] $end
$var wire 1 HA l2_2_s [32] $end
$var wire 1 IA l2_2_s [31] $end
$var wire 1 JA l2_2_s [30] $end
$var wire 1 KA l2_2_s [29] $end
$var wire 1 LA l2_2_s [28] $end
$var wire 1 MA l2_2_s [27] $end
$var wire 1 NA l2_2_s [26] $end
$var wire 1 OA l2_2_s [25] $end
$var wire 1 PA l2_2_s [24] $end
$var wire 1 QA l2_2_s [23] $end
$var wire 1 RA l2_2_s [22] $end
$var wire 1 SA l2_2_s [21] $end
$var wire 1 TA l2_2_s [20] $end
$var wire 1 UA l2_2_s [19] $end
$var wire 1 VA l2_2_s [18] $end
$var wire 1 WA l2_2_s [17] $end
$var wire 1 XA l2_2_s [16] $end
$var wire 1 YA l2_2_s [15] $end
$var wire 1 ZA l2_2_s [14] $end
$var wire 1 [A l2_2_s [13] $end
$var wire 1 \A l2_2_s [12] $end
$var wire 1 ]A l2_2_s [11] $end
$var wire 1 ^A l2_2_s [10] $end
$var wire 1 _A l2_2_s [9] $end
$var wire 1 `A l2_2_s [8] $end
$var wire 1 aA l2_2_s [7] $end
$var wire 1 bA l2_2_s [6] $end
$var wire 1 cA l2_2_s [5] $end
$var wire 1 dA l2_2_s [4] $end
$var wire 1 eA l2_2_s [3] $end
$var wire 1 fA l2_2_s [2] $end
$var wire 1 gA l2_2_s [1] $end
$var wire 1 hA l2_2_s [0] $end
$var wire 1 iA l2_2_ca [46] $end
$var wire 1 jA l2_2_ca [45] $end
$var wire 1 kA l2_2_ca [44] $end
$var wire 1 lA l2_2_ca [43] $end
$var wire 1 mA l2_2_ca [42] $end
$var wire 1 nA l2_2_ca [41] $end
$var wire 1 oA l2_2_ca [40] $end
$var wire 1 pA l2_2_ca [39] $end
$var wire 1 qA l2_2_ca [38] $end
$var wire 1 rA l2_2_ca [37] $end
$var wire 1 sA l2_2_ca [36] $end
$var wire 1 tA l2_2_ca [35] $end
$var wire 1 uA l2_2_ca [34] $end
$var wire 1 vA l2_2_ca [33] $end
$var wire 1 wA l2_2_ca [32] $end
$var wire 1 xA l2_2_ca [31] $end
$var wire 1 yA l2_2_ca [30] $end
$var wire 1 zA l2_2_ca [29] $end
$var wire 1 {A l2_2_ca [28] $end
$var wire 1 |A l2_2_ca [27] $end
$var wire 1 }A l2_2_ca [26] $end
$var wire 1 ~A l2_2_ca [25] $end
$var wire 1 !B l2_2_ca [24] $end
$var wire 1 "B l2_2_ca [23] $end
$var wire 1 #B l2_2_ca [22] $end
$var wire 1 $B l2_2_ca [21] $end
$var wire 1 %B l2_2_ca [20] $end
$var wire 1 &B l2_2_ca [19] $end
$var wire 1 'B l2_2_ca [18] $end
$var wire 1 (B l2_2_ca [17] $end
$var wire 1 )B l2_2_ca [16] $end
$var wire 1 *B l2_2_ca [15] $end
$var wire 1 +B l2_2_ca [14] $end
$var wire 1 ,B l2_2_ca [13] $end
$var wire 1 -B l2_2_ca [12] $end
$var wire 1 .B l2_2_ca [11] $end
$var wire 1 /B l2_2_ca [10] $end
$var wire 1 0B l2_2_ca [9] $end
$var wire 1 1B l2_2_ca [8] $end
$var wire 1 2B l2_2_ca [7] $end
$var wire 1 3B l2_2_ca [6] $end
$var wire 1 4B l2_2_ca [5] $end
$var wire 1 5B l2_2_ca [4] $end
$var wire 1 6B l2_2_ca [3] $end
$var wire 1 7B l2_2_ca [2] $end
$var wire 1 8B l2_2_ca [1] $end
$var wire 1 9B l2_2_ca [0] $end
$var wire 1 :B l2_3_0 [43] $end
$var wire 1 ;B l2_3_0 [42] $end
$var wire 1 <B l2_3_0 [41] $end
$var wire 1 =B l2_3_0 [40] $end
$var wire 1 >B l2_3_0 [39] $end
$var wire 1 ?B l2_3_0 [38] $end
$var wire 1 @B l2_3_0 [37] $end
$var wire 1 AB l2_3_0 [36] $end
$var wire 1 BB l2_3_0 [35] $end
$var wire 1 CB l2_3_0 [34] $end
$var wire 1 DB l2_3_0 [33] $end
$var wire 1 EB l2_3_0 [32] $end
$var wire 1 FB l2_3_0 [31] $end
$var wire 1 GB l2_3_0 [30] $end
$var wire 1 HB l2_3_0 [29] $end
$var wire 1 IB l2_3_0 [28] $end
$var wire 1 JB l2_3_0 [27] $end
$var wire 1 KB l2_3_0 [26] $end
$var wire 1 LB l2_3_0 [25] $end
$var wire 1 MB l2_3_0 [24] $end
$var wire 1 NB l2_3_0 [23] $end
$var wire 1 OB l2_3_0 [22] $end
$var wire 1 PB l2_3_0 [21] $end
$var wire 1 QB l2_3_0 [20] $end
$var wire 1 RB l2_3_0 [19] $end
$var wire 1 SB l2_3_0 [18] $end
$var wire 1 TB l2_3_0 [17] $end
$var wire 1 UB l2_3_0 [16] $end
$var wire 1 VB l2_3_0 [15] $end
$var wire 1 WB l2_3_0 [14] $end
$var wire 1 XB l2_3_0 [13] $end
$var wire 1 YB l2_3_0 [12] $end
$var wire 1 ZB l2_3_0 [11] $end
$var wire 1 [B l2_3_0 [10] $end
$var wire 1 \B l2_3_0 [9] $end
$var wire 1 ]B l2_3_0 [8] $end
$var wire 1 ^B l2_3_0 [7] $end
$var wire 1 _B l2_3_0 [6] $end
$var wire 1 `B l2_3_0 [5] $end
$var wire 1 aB l2_3_0 [4] $end
$var wire 1 bB l2_3_0 [3] $end
$var wire 1 cB l2_3_0 [2] $end
$var wire 1 dB l2_3_0 [1] $end
$var wire 1 eB l2_3_0 [0] $end
$var wire 1 fB l2_3_1 [43] $end
$var wire 1 gB l2_3_1 [42] $end
$var wire 1 hB l2_3_1 [41] $end
$var wire 1 iB l2_3_1 [40] $end
$var wire 1 jB l2_3_1 [39] $end
$var wire 1 kB l2_3_1 [38] $end
$var wire 1 lB l2_3_1 [37] $end
$var wire 1 mB l2_3_1 [36] $end
$var wire 1 nB l2_3_1 [35] $end
$var wire 1 oB l2_3_1 [34] $end
$var wire 1 pB l2_3_1 [33] $end
$var wire 1 qB l2_3_1 [32] $end
$var wire 1 rB l2_3_1 [31] $end
$var wire 1 sB l2_3_1 [30] $end
$var wire 1 tB l2_3_1 [29] $end
$var wire 1 uB l2_3_1 [28] $end
$var wire 1 vB l2_3_1 [27] $end
$var wire 1 wB l2_3_1 [26] $end
$var wire 1 xB l2_3_1 [25] $end
$var wire 1 yB l2_3_1 [24] $end
$var wire 1 zB l2_3_1 [23] $end
$var wire 1 {B l2_3_1 [22] $end
$var wire 1 |B l2_3_1 [21] $end
$var wire 1 }B l2_3_1 [20] $end
$var wire 1 ~B l2_3_1 [19] $end
$var wire 1 !C l2_3_1 [18] $end
$var wire 1 "C l2_3_1 [17] $end
$var wire 1 #C l2_3_1 [16] $end
$var wire 1 $C l2_3_1 [15] $end
$var wire 1 %C l2_3_1 [14] $end
$var wire 1 &C l2_3_1 [13] $end
$var wire 1 'C l2_3_1 [12] $end
$var wire 1 (C l2_3_1 [11] $end
$var wire 1 )C l2_3_1 [10] $end
$var wire 1 *C l2_3_1 [9] $end
$var wire 1 +C l2_3_1 [8] $end
$var wire 1 ,C l2_3_1 [7] $end
$var wire 1 -C l2_3_1 [6] $end
$var wire 1 .C l2_3_1 [5] $end
$var wire 1 /C l2_3_1 [4] $end
$var wire 1 0C l2_3_1 [3] $end
$var wire 1 1C l2_3_1 [2] $end
$var wire 1 2C l2_3_1 [1] $end
$var wire 1 3C l2_3_1 [0] $end
$var wire 1 4C l2_3_2 [43] $end
$var wire 1 5C l2_3_2 [42] $end
$var wire 1 6C l2_3_2 [41] $end
$var wire 1 7C l2_3_2 [40] $end
$var wire 1 8C l2_3_2 [39] $end
$var wire 1 9C l2_3_2 [38] $end
$var wire 1 :C l2_3_2 [37] $end
$var wire 1 ;C l2_3_2 [36] $end
$var wire 1 <C l2_3_2 [35] $end
$var wire 1 =C l2_3_2 [34] $end
$var wire 1 >C l2_3_2 [33] $end
$var wire 1 ?C l2_3_2 [32] $end
$var wire 1 @C l2_3_2 [31] $end
$var wire 1 AC l2_3_2 [30] $end
$var wire 1 BC l2_3_2 [29] $end
$var wire 1 CC l2_3_2 [28] $end
$var wire 1 DC l2_3_2 [27] $end
$var wire 1 EC l2_3_2 [26] $end
$var wire 1 FC l2_3_2 [25] $end
$var wire 1 GC l2_3_2 [24] $end
$var wire 1 HC l2_3_2 [23] $end
$var wire 1 IC l2_3_2 [22] $end
$var wire 1 JC l2_3_2 [21] $end
$var wire 1 KC l2_3_2 [20] $end
$var wire 1 LC l2_3_2 [19] $end
$var wire 1 MC l2_3_2 [18] $end
$var wire 1 NC l2_3_2 [17] $end
$var wire 1 OC l2_3_2 [16] $end
$var wire 1 PC l2_3_2 [15] $end
$var wire 1 QC l2_3_2 [14] $end
$var wire 1 RC l2_3_2 [13] $end
$var wire 1 SC l2_3_2 [12] $end
$var wire 1 TC l2_3_2 [11] $end
$var wire 1 UC l2_3_2 [10] $end
$var wire 1 VC l2_3_2 [9] $end
$var wire 1 WC l2_3_2 [8] $end
$var wire 1 XC l2_3_2 [7] $end
$var wire 1 YC l2_3_2 [6] $end
$var wire 1 ZC l2_3_2 [5] $end
$var wire 1 [C l2_3_2 [4] $end
$var wire 1 \C l2_3_2 [3] $end
$var wire 1 ]C l2_3_2 [2] $end
$var wire 1 ^C l2_3_2 [1] $end
$var wire 1 _C l2_3_2 [0] $end
$var wire 1 `C l2_3_3 [43] $end
$var wire 1 aC l2_3_3 [42] $end
$var wire 1 bC l2_3_3 [41] $end
$var wire 1 cC l2_3_3 [40] $end
$var wire 1 dC l2_3_3 [39] $end
$var wire 1 eC l2_3_3 [38] $end
$var wire 1 fC l2_3_3 [37] $end
$var wire 1 gC l2_3_3 [36] $end
$var wire 1 hC l2_3_3 [35] $end
$var wire 1 iC l2_3_3 [34] $end
$var wire 1 jC l2_3_3 [33] $end
$var wire 1 kC l2_3_3 [32] $end
$var wire 1 lC l2_3_3 [31] $end
$var wire 1 mC l2_3_3 [30] $end
$var wire 1 nC l2_3_3 [29] $end
$var wire 1 oC l2_3_3 [28] $end
$var wire 1 pC l2_3_3 [27] $end
$var wire 1 qC l2_3_3 [26] $end
$var wire 1 rC l2_3_3 [25] $end
$var wire 1 sC l2_3_3 [24] $end
$var wire 1 tC l2_3_3 [23] $end
$var wire 1 uC l2_3_3 [22] $end
$var wire 1 vC l2_3_3 [21] $end
$var wire 1 wC l2_3_3 [20] $end
$var wire 1 xC l2_3_3 [19] $end
$var wire 1 yC l2_3_3 [18] $end
$var wire 1 zC l2_3_3 [17] $end
$var wire 1 {C l2_3_3 [16] $end
$var wire 1 |C l2_3_3 [15] $end
$var wire 1 }C l2_3_3 [14] $end
$var wire 1 ~C l2_3_3 [13] $end
$var wire 1 !D l2_3_3 [12] $end
$var wire 1 "D l2_3_3 [11] $end
$var wire 1 #D l2_3_3 [10] $end
$var wire 1 $D l2_3_3 [9] $end
$var wire 1 %D l2_3_3 [8] $end
$var wire 1 &D l2_3_3 [7] $end
$var wire 1 'D l2_3_3 [6] $end
$var wire 1 (D l2_3_3 [5] $end
$var wire 1 )D l2_3_3 [4] $end
$var wire 1 *D l2_3_3 [3] $end
$var wire 1 +D l2_3_3 [2] $end
$var wire 1 ,D l2_3_3 [1] $end
$var wire 1 -D l2_3_3 [0] $end
$var wire 1 .D l2_3_cin [43] $end
$var wire 1 /D l2_3_cin [42] $end
$var wire 1 0D l2_3_cin [41] $end
$var wire 1 1D l2_3_cin [40] $end
$var wire 1 2D l2_3_cin [39] $end
$var wire 1 3D l2_3_cin [38] $end
$var wire 1 4D l2_3_cin [37] $end
$var wire 1 5D l2_3_cin [36] $end
$var wire 1 6D l2_3_cin [35] $end
$var wire 1 7D l2_3_cin [34] $end
$var wire 1 8D l2_3_cin [33] $end
$var wire 1 9D l2_3_cin [32] $end
$var wire 1 :D l2_3_cin [31] $end
$var wire 1 ;D l2_3_cin [30] $end
$var wire 1 <D l2_3_cin [29] $end
$var wire 1 =D l2_3_cin [28] $end
$var wire 1 >D l2_3_cin [27] $end
$var wire 1 ?D l2_3_cin [26] $end
$var wire 1 @D l2_3_cin [25] $end
$var wire 1 AD l2_3_cin [24] $end
$var wire 1 BD l2_3_cin [23] $end
$var wire 1 CD l2_3_cin [22] $end
$var wire 1 DD l2_3_cin [21] $end
$var wire 1 ED l2_3_cin [20] $end
$var wire 1 FD l2_3_cin [19] $end
$var wire 1 GD l2_3_cin [18] $end
$var wire 1 HD l2_3_cin [17] $end
$var wire 1 ID l2_3_cin [16] $end
$var wire 1 JD l2_3_cin [15] $end
$var wire 1 KD l2_3_cin [14] $end
$var wire 1 LD l2_3_cin [13] $end
$var wire 1 MD l2_3_cin [12] $end
$var wire 1 ND l2_3_cin [11] $end
$var wire 1 OD l2_3_cin [10] $end
$var wire 1 PD l2_3_cin [9] $end
$var wire 1 QD l2_3_cin [8] $end
$var wire 1 RD l2_3_cin [7] $end
$var wire 1 SD l2_3_cin [6] $end
$var wire 1 TD l2_3_cin [5] $end
$var wire 1 UD l2_3_cin [4] $end
$var wire 1 VD l2_3_cin [3] $end
$var wire 1 WD l2_3_cin [2] $end
$var wire 1 XD l2_3_cin [1] $end
$var wire 1 YD l2_3_cin [0] $end
$var wire 1 ZD l2_3_cout [43] $end
$var wire 1 [D l2_3_cout [42] $end
$var wire 1 \D l2_3_cout [41] $end
$var wire 1 ]D l2_3_cout [40] $end
$var wire 1 ^D l2_3_cout [39] $end
$var wire 1 _D l2_3_cout [38] $end
$var wire 1 `D l2_3_cout [37] $end
$var wire 1 aD l2_3_cout [36] $end
$var wire 1 bD l2_3_cout [35] $end
$var wire 1 cD l2_3_cout [34] $end
$var wire 1 dD l2_3_cout [33] $end
$var wire 1 eD l2_3_cout [32] $end
$var wire 1 fD l2_3_cout [31] $end
$var wire 1 gD l2_3_cout [30] $end
$var wire 1 hD l2_3_cout [29] $end
$var wire 1 iD l2_3_cout [28] $end
$var wire 1 jD l2_3_cout [27] $end
$var wire 1 kD l2_3_cout [26] $end
$var wire 1 lD l2_3_cout [25] $end
$var wire 1 mD l2_3_cout [24] $end
$var wire 1 nD l2_3_cout [23] $end
$var wire 1 oD l2_3_cout [22] $end
$var wire 1 pD l2_3_cout [21] $end
$var wire 1 qD l2_3_cout [20] $end
$var wire 1 rD l2_3_cout [19] $end
$var wire 1 sD l2_3_cout [18] $end
$var wire 1 tD l2_3_cout [17] $end
$var wire 1 uD l2_3_cout [16] $end
$var wire 1 vD l2_3_cout [15] $end
$var wire 1 wD l2_3_cout [14] $end
$var wire 1 xD l2_3_cout [13] $end
$var wire 1 yD l2_3_cout [12] $end
$var wire 1 zD l2_3_cout [11] $end
$var wire 1 {D l2_3_cout [10] $end
$var wire 1 |D l2_3_cout [9] $end
$var wire 1 }D l2_3_cout [8] $end
$var wire 1 ~D l2_3_cout [7] $end
$var wire 1 !E l2_3_cout [6] $end
$var wire 1 "E l2_3_cout [5] $end
$var wire 1 #E l2_3_cout [4] $end
$var wire 1 $E l2_3_cout [3] $end
$var wire 1 %E l2_3_cout [2] $end
$var wire 1 &E l2_3_cout [1] $end
$var wire 1 'E l2_3_cout [0] $end
$var wire 1 (E l2_3_s [43] $end
$var wire 1 )E l2_3_s [42] $end
$var wire 1 *E l2_3_s [41] $end
$var wire 1 +E l2_3_s [40] $end
$var wire 1 ,E l2_3_s [39] $end
$var wire 1 -E l2_3_s [38] $end
$var wire 1 .E l2_3_s [37] $end
$var wire 1 /E l2_3_s [36] $end
$var wire 1 0E l2_3_s [35] $end
$var wire 1 1E l2_3_s [34] $end
$var wire 1 2E l2_3_s [33] $end
$var wire 1 3E l2_3_s [32] $end
$var wire 1 4E l2_3_s [31] $end
$var wire 1 5E l2_3_s [30] $end
$var wire 1 6E l2_3_s [29] $end
$var wire 1 7E l2_3_s [28] $end
$var wire 1 8E l2_3_s [27] $end
$var wire 1 9E l2_3_s [26] $end
$var wire 1 :E l2_3_s [25] $end
$var wire 1 ;E l2_3_s [24] $end
$var wire 1 <E l2_3_s [23] $end
$var wire 1 =E l2_3_s [22] $end
$var wire 1 >E l2_3_s [21] $end
$var wire 1 ?E l2_3_s [20] $end
$var wire 1 @E l2_3_s [19] $end
$var wire 1 AE l2_3_s [18] $end
$var wire 1 BE l2_3_s [17] $end
$var wire 1 CE l2_3_s [16] $end
$var wire 1 DE l2_3_s [15] $end
$var wire 1 EE l2_3_s [14] $end
$var wire 1 FE l2_3_s [13] $end
$var wire 1 GE l2_3_s [12] $end
$var wire 1 HE l2_3_s [11] $end
$var wire 1 IE l2_3_s [10] $end
$var wire 1 JE l2_3_s [9] $end
$var wire 1 KE l2_3_s [8] $end
$var wire 1 LE l2_3_s [7] $end
$var wire 1 ME l2_3_s [6] $end
$var wire 1 NE l2_3_s [5] $end
$var wire 1 OE l2_3_s [4] $end
$var wire 1 PE l2_3_s [3] $end
$var wire 1 QE l2_3_s [2] $end
$var wire 1 RE l2_3_s [1] $end
$var wire 1 SE l2_3_s [0] $end
$var wire 1 TE l2_3_ca [43] $end
$var wire 1 UE l2_3_ca [42] $end
$var wire 1 VE l2_3_ca [41] $end
$var wire 1 WE l2_3_ca [40] $end
$var wire 1 XE l2_3_ca [39] $end
$var wire 1 YE l2_3_ca [38] $end
$var wire 1 ZE l2_3_ca [37] $end
$var wire 1 [E l2_3_ca [36] $end
$var wire 1 \E l2_3_ca [35] $end
$var wire 1 ]E l2_3_ca [34] $end
$var wire 1 ^E l2_3_ca [33] $end
$var wire 1 _E l2_3_ca [32] $end
$var wire 1 `E l2_3_ca [31] $end
$var wire 1 aE l2_3_ca [30] $end
$var wire 1 bE l2_3_ca [29] $end
$var wire 1 cE l2_3_ca [28] $end
$var wire 1 dE l2_3_ca [27] $end
$var wire 1 eE l2_3_ca [26] $end
$var wire 1 fE l2_3_ca [25] $end
$var wire 1 gE l2_3_ca [24] $end
$var wire 1 hE l2_3_ca [23] $end
$var wire 1 iE l2_3_ca [22] $end
$var wire 1 jE l2_3_ca [21] $end
$var wire 1 kE l2_3_ca [20] $end
$var wire 1 lE l2_3_ca [19] $end
$var wire 1 mE l2_3_ca [18] $end
$var wire 1 nE l2_3_ca [17] $end
$var wire 1 oE l2_3_ca [16] $end
$var wire 1 pE l2_3_ca [15] $end
$var wire 1 qE l2_3_ca [14] $end
$var wire 1 rE l2_3_ca [13] $end
$var wire 1 sE l2_3_ca [12] $end
$var wire 1 tE l2_3_ca [11] $end
$var wire 1 uE l2_3_ca [10] $end
$var wire 1 vE l2_3_ca [9] $end
$var wire 1 wE l2_3_ca [8] $end
$var wire 1 xE l2_3_ca [7] $end
$var wire 1 yE l2_3_ca [6] $end
$var wire 1 zE l2_3_ca [5] $end
$var wire 1 {E l2_3_ca [4] $end
$var wire 1 |E l2_3_ca [3] $end
$var wire 1 }E l2_3_ca [2] $end
$var wire 1 ~E l2_3_ca [1] $end
$var wire 1 !F l2_3_ca [0] $end
$var reg 43 "F l2_s1_reg [42:0] $end
$var reg 43 #F l2_c1_reg [42:0] $end
$var reg 47 $F l2_s2_reg [46:0] $end
$var reg 47 %F l2_c2_reg [46:0] $end
$var reg 44 &F l2_s3_reg [43:0] $end
$var reg 44 'F l2_c3_reg [43:0] $end
$var wire 1 (F l3_1_0 [54] $end
$var wire 1 )F l3_1_0 [53] $end
$var wire 1 *F l3_1_0 [52] $end
$var wire 1 +F l3_1_0 [51] $end
$var wire 1 ,F l3_1_0 [50] $end
$var wire 1 -F l3_1_0 [49] $end
$var wire 1 .F l3_1_0 [48] $end
$var wire 1 /F l3_1_0 [47] $end
$var wire 1 0F l3_1_0 [46] $end
$var wire 1 1F l3_1_0 [45] $end
$var wire 1 2F l3_1_0 [44] $end
$var wire 1 3F l3_1_0 [43] $end
$var wire 1 4F l3_1_0 [42] $end
$var wire 1 5F l3_1_0 [41] $end
$var wire 1 6F l3_1_0 [40] $end
$var wire 1 7F l3_1_0 [39] $end
$var wire 1 8F l3_1_0 [38] $end
$var wire 1 9F l3_1_0 [37] $end
$var wire 1 :F l3_1_0 [36] $end
$var wire 1 ;F l3_1_0 [35] $end
$var wire 1 <F l3_1_0 [34] $end
$var wire 1 =F l3_1_0 [33] $end
$var wire 1 >F l3_1_0 [32] $end
$var wire 1 ?F l3_1_0 [31] $end
$var wire 1 @F l3_1_0 [30] $end
$var wire 1 AF l3_1_0 [29] $end
$var wire 1 BF l3_1_0 [28] $end
$var wire 1 CF l3_1_0 [27] $end
$var wire 1 DF l3_1_0 [26] $end
$var wire 1 EF l3_1_0 [25] $end
$var wire 1 FF l3_1_0 [24] $end
$var wire 1 GF l3_1_0 [23] $end
$var wire 1 HF l3_1_0 [22] $end
$var wire 1 IF l3_1_0 [21] $end
$var wire 1 JF l3_1_0 [20] $end
$var wire 1 KF l3_1_0 [19] $end
$var wire 1 LF l3_1_0 [18] $end
$var wire 1 MF l3_1_0 [17] $end
$var wire 1 NF l3_1_0 [16] $end
$var wire 1 OF l3_1_0 [15] $end
$var wire 1 PF l3_1_0 [14] $end
$var wire 1 QF l3_1_0 [13] $end
$var wire 1 RF l3_1_0 [12] $end
$var wire 1 SF l3_1_0 [11] $end
$var wire 1 TF l3_1_0 [10] $end
$var wire 1 UF l3_1_0 [9] $end
$var wire 1 VF l3_1_0 [8] $end
$var wire 1 WF l3_1_0 [7] $end
$var wire 1 XF l3_1_0 [6] $end
$var wire 1 YF l3_1_0 [5] $end
$var wire 1 ZF l3_1_0 [4] $end
$var wire 1 [F l3_1_0 [3] $end
$var wire 1 \F l3_1_0 [2] $end
$var wire 1 ]F l3_1_0 [1] $end
$var wire 1 ^F l3_1_0 [0] $end
$var wire 1 _F l3_1_1 [54] $end
$var wire 1 `F l3_1_1 [53] $end
$var wire 1 aF l3_1_1 [52] $end
$var wire 1 bF l3_1_1 [51] $end
$var wire 1 cF l3_1_1 [50] $end
$var wire 1 dF l3_1_1 [49] $end
$var wire 1 eF l3_1_1 [48] $end
$var wire 1 fF l3_1_1 [47] $end
$var wire 1 gF l3_1_1 [46] $end
$var wire 1 hF l3_1_1 [45] $end
$var wire 1 iF l3_1_1 [44] $end
$var wire 1 jF l3_1_1 [43] $end
$var wire 1 kF l3_1_1 [42] $end
$var wire 1 lF l3_1_1 [41] $end
$var wire 1 mF l3_1_1 [40] $end
$var wire 1 nF l3_1_1 [39] $end
$var wire 1 oF l3_1_1 [38] $end
$var wire 1 pF l3_1_1 [37] $end
$var wire 1 qF l3_1_1 [36] $end
$var wire 1 rF l3_1_1 [35] $end
$var wire 1 sF l3_1_1 [34] $end
$var wire 1 tF l3_1_1 [33] $end
$var wire 1 uF l3_1_1 [32] $end
$var wire 1 vF l3_1_1 [31] $end
$var wire 1 wF l3_1_1 [30] $end
$var wire 1 xF l3_1_1 [29] $end
$var wire 1 yF l3_1_1 [28] $end
$var wire 1 zF l3_1_1 [27] $end
$var wire 1 {F l3_1_1 [26] $end
$var wire 1 |F l3_1_1 [25] $end
$var wire 1 }F l3_1_1 [24] $end
$var wire 1 ~F l3_1_1 [23] $end
$var wire 1 !G l3_1_1 [22] $end
$var wire 1 "G l3_1_1 [21] $end
$var wire 1 #G l3_1_1 [20] $end
$var wire 1 $G l3_1_1 [19] $end
$var wire 1 %G l3_1_1 [18] $end
$var wire 1 &G l3_1_1 [17] $end
$var wire 1 'G l3_1_1 [16] $end
$var wire 1 (G l3_1_1 [15] $end
$var wire 1 )G l3_1_1 [14] $end
$var wire 1 *G l3_1_1 [13] $end
$var wire 1 +G l3_1_1 [12] $end
$var wire 1 ,G l3_1_1 [11] $end
$var wire 1 -G l3_1_1 [10] $end
$var wire 1 .G l3_1_1 [9] $end
$var wire 1 /G l3_1_1 [8] $end
$var wire 1 0G l3_1_1 [7] $end
$var wire 1 1G l3_1_1 [6] $end
$var wire 1 2G l3_1_1 [5] $end
$var wire 1 3G l3_1_1 [4] $end
$var wire 1 4G l3_1_1 [3] $end
$var wire 1 5G l3_1_1 [2] $end
$var wire 1 6G l3_1_1 [1] $end
$var wire 1 7G l3_1_1 [0] $end
$var wire 1 8G l3_1_2 [54] $end
$var wire 1 9G l3_1_2 [53] $end
$var wire 1 :G l3_1_2 [52] $end
$var wire 1 ;G l3_1_2 [51] $end
$var wire 1 <G l3_1_2 [50] $end
$var wire 1 =G l3_1_2 [49] $end
$var wire 1 >G l3_1_2 [48] $end
$var wire 1 ?G l3_1_2 [47] $end
$var wire 1 @G l3_1_2 [46] $end
$var wire 1 AG l3_1_2 [45] $end
$var wire 1 BG l3_1_2 [44] $end
$var wire 1 CG l3_1_2 [43] $end
$var wire 1 DG l3_1_2 [42] $end
$var wire 1 EG l3_1_2 [41] $end
$var wire 1 FG l3_1_2 [40] $end
$var wire 1 GG l3_1_2 [39] $end
$var wire 1 HG l3_1_2 [38] $end
$var wire 1 IG l3_1_2 [37] $end
$var wire 1 JG l3_1_2 [36] $end
$var wire 1 KG l3_1_2 [35] $end
$var wire 1 LG l3_1_2 [34] $end
$var wire 1 MG l3_1_2 [33] $end
$var wire 1 NG l3_1_2 [32] $end
$var wire 1 OG l3_1_2 [31] $end
$var wire 1 PG l3_1_2 [30] $end
$var wire 1 QG l3_1_2 [29] $end
$var wire 1 RG l3_1_2 [28] $end
$var wire 1 SG l3_1_2 [27] $end
$var wire 1 TG l3_1_2 [26] $end
$var wire 1 UG l3_1_2 [25] $end
$var wire 1 VG l3_1_2 [24] $end
$var wire 1 WG l3_1_2 [23] $end
$var wire 1 XG l3_1_2 [22] $end
$var wire 1 YG l3_1_2 [21] $end
$var wire 1 ZG l3_1_2 [20] $end
$var wire 1 [G l3_1_2 [19] $end
$var wire 1 \G l3_1_2 [18] $end
$var wire 1 ]G l3_1_2 [17] $end
$var wire 1 ^G l3_1_2 [16] $end
$var wire 1 _G l3_1_2 [15] $end
$var wire 1 `G l3_1_2 [14] $end
$var wire 1 aG l3_1_2 [13] $end
$var wire 1 bG l3_1_2 [12] $end
$var wire 1 cG l3_1_2 [11] $end
$var wire 1 dG l3_1_2 [10] $end
$var wire 1 eG l3_1_2 [9] $end
$var wire 1 fG l3_1_2 [8] $end
$var wire 1 gG l3_1_2 [7] $end
$var wire 1 hG l3_1_2 [6] $end
$var wire 1 iG l3_1_2 [5] $end
$var wire 1 jG l3_1_2 [4] $end
$var wire 1 kG l3_1_2 [3] $end
$var wire 1 lG l3_1_2 [2] $end
$var wire 1 mG l3_1_2 [1] $end
$var wire 1 nG l3_1_2 [0] $end
$var wire 1 oG l3_1_s [54] $end
$var wire 1 pG l3_1_s [53] $end
$var wire 1 qG l3_1_s [52] $end
$var wire 1 rG l3_1_s [51] $end
$var wire 1 sG l3_1_s [50] $end
$var wire 1 tG l3_1_s [49] $end
$var wire 1 uG l3_1_s [48] $end
$var wire 1 vG l3_1_s [47] $end
$var wire 1 wG l3_1_s [46] $end
$var wire 1 xG l3_1_s [45] $end
$var wire 1 yG l3_1_s [44] $end
$var wire 1 zG l3_1_s [43] $end
$var wire 1 {G l3_1_s [42] $end
$var wire 1 |G l3_1_s [41] $end
$var wire 1 }G l3_1_s [40] $end
$var wire 1 ~G l3_1_s [39] $end
$var wire 1 !H l3_1_s [38] $end
$var wire 1 "H l3_1_s [37] $end
$var wire 1 #H l3_1_s [36] $end
$var wire 1 $H l3_1_s [35] $end
$var wire 1 %H l3_1_s [34] $end
$var wire 1 &H l3_1_s [33] $end
$var wire 1 'H l3_1_s [32] $end
$var wire 1 (H l3_1_s [31] $end
$var wire 1 )H l3_1_s [30] $end
$var wire 1 *H l3_1_s [29] $end
$var wire 1 +H l3_1_s [28] $end
$var wire 1 ,H l3_1_s [27] $end
$var wire 1 -H l3_1_s [26] $end
$var wire 1 .H l3_1_s [25] $end
$var wire 1 /H l3_1_s [24] $end
$var wire 1 0H l3_1_s [23] $end
$var wire 1 1H l3_1_s [22] $end
$var wire 1 2H l3_1_s [21] $end
$var wire 1 3H l3_1_s [20] $end
$var wire 1 4H l3_1_s [19] $end
$var wire 1 5H l3_1_s [18] $end
$var wire 1 6H l3_1_s [17] $end
$var wire 1 7H l3_1_s [16] $end
$var wire 1 8H l3_1_s [15] $end
$var wire 1 9H l3_1_s [14] $end
$var wire 1 :H l3_1_s [13] $end
$var wire 1 ;H l3_1_s [12] $end
$var wire 1 <H l3_1_s [11] $end
$var wire 1 =H l3_1_s [10] $end
$var wire 1 >H l3_1_s [9] $end
$var wire 1 ?H l3_1_s [8] $end
$var wire 1 @H l3_1_s [7] $end
$var wire 1 AH l3_1_s [6] $end
$var wire 1 BH l3_1_s [5] $end
$var wire 1 CH l3_1_s [4] $end
$var wire 1 DH l3_1_s [3] $end
$var wire 1 EH l3_1_s [2] $end
$var wire 1 FH l3_1_s [1] $end
$var wire 1 GH l3_1_s [0] $end
$var wire 1 HH l3_1_ca [54] $end
$var wire 1 IH l3_1_ca [53] $end
$var wire 1 JH l3_1_ca [52] $end
$var wire 1 KH l3_1_ca [51] $end
$var wire 1 LH l3_1_ca [50] $end
$var wire 1 MH l3_1_ca [49] $end
$var wire 1 NH l3_1_ca [48] $end
$var wire 1 OH l3_1_ca [47] $end
$var wire 1 PH l3_1_ca [46] $end
$var wire 1 QH l3_1_ca [45] $end
$var wire 1 RH l3_1_ca [44] $end
$var wire 1 SH l3_1_ca [43] $end
$var wire 1 TH l3_1_ca [42] $end
$var wire 1 UH l3_1_ca [41] $end
$var wire 1 VH l3_1_ca [40] $end
$var wire 1 WH l3_1_ca [39] $end
$var wire 1 XH l3_1_ca [38] $end
$var wire 1 YH l3_1_ca [37] $end
$var wire 1 ZH l3_1_ca [36] $end
$var wire 1 [H l3_1_ca [35] $end
$var wire 1 \H l3_1_ca [34] $end
$var wire 1 ]H l3_1_ca [33] $end
$var wire 1 ^H l3_1_ca [32] $end
$var wire 1 _H l3_1_ca [31] $end
$var wire 1 `H l3_1_ca [30] $end
$var wire 1 aH l3_1_ca [29] $end
$var wire 1 bH l3_1_ca [28] $end
$var wire 1 cH l3_1_ca [27] $end
$var wire 1 dH l3_1_ca [26] $end
$var wire 1 eH l3_1_ca [25] $end
$var wire 1 fH l3_1_ca [24] $end
$var wire 1 gH l3_1_ca [23] $end
$var wire 1 hH l3_1_ca [22] $end
$var wire 1 iH l3_1_ca [21] $end
$var wire 1 jH l3_1_ca [20] $end
$var wire 1 kH l3_1_ca [19] $end
$var wire 1 lH l3_1_ca [18] $end
$var wire 1 mH l3_1_ca [17] $end
$var wire 1 nH l3_1_ca [16] $end
$var wire 1 oH l3_1_ca [15] $end
$var wire 1 pH l3_1_ca [14] $end
$var wire 1 qH l3_1_ca [13] $end
$var wire 1 rH l3_1_ca [12] $end
$var wire 1 sH l3_1_ca [11] $end
$var wire 1 tH l3_1_ca [10] $end
$var wire 1 uH l3_1_ca [9] $end
$var wire 1 vH l3_1_ca [8] $end
$var wire 1 wH l3_1_ca [7] $end
$var wire 1 xH l3_1_ca [6] $end
$var wire 1 yH l3_1_ca [5] $end
$var wire 1 zH l3_1_ca [4] $end
$var wire 1 {H l3_1_ca [3] $end
$var wire 1 |H l3_1_ca [2] $end
$var wire 1 }H l3_1_ca [1] $end
$var wire 1 ~H l3_1_ca [0] $end
$var wire 1 !I l3_2_0 [54] $end
$var wire 1 "I l3_2_0 [53] $end
$var wire 1 #I l3_2_0 [52] $end
$var wire 1 $I l3_2_0 [51] $end
$var wire 1 %I l3_2_0 [50] $end
$var wire 1 &I l3_2_0 [49] $end
$var wire 1 'I l3_2_0 [48] $end
$var wire 1 (I l3_2_0 [47] $end
$var wire 1 )I l3_2_0 [46] $end
$var wire 1 *I l3_2_0 [45] $end
$var wire 1 +I l3_2_0 [44] $end
$var wire 1 ,I l3_2_0 [43] $end
$var wire 1 -I l3_2_0 [42] $end
$var wire 1 .I l3_2_0 [41] $end
$var wire 1 /I l3_2_0 [40] $end
$var wire 1 0I l3_2_0 [39] $end
$var wire 1 1I l3_2_0 [38] $end
$var wire 1 2I l3_2_0 [37] $end
$var wire 1 3I l3_2_0 [36] $end
$var wire 1 4I l3_2_0 [35] $end
$var wire 1 5I l3_2_0 [34] $end
$var wire 1 6I l3_2_0 [33] $end
$var wire 1 7I l3_2_0 [32] $end
$var wire 1 8I l3_2_0 [31] $end
$var wire 1 9I l3_2_0 [30] $end
$var wire 1 :I l3_2_0 [29] $end
$var wire 1 ;I l3_2_0 [28] $end
$var wire 1 <I l3_2_0 [27] $end
$var wire 1 =I l3_2_0 [26] $end
$var wire 1 >I l3_2_0 [25] $end
$var wire 1 ?I l3_2_0 [24] $end
$var wire 1 @I l3_2_0 [23] $end
$var wire 1 AI l3_2_0 [22] $end
$var wire 1 BI l3_2_0 [21] $end
$var wire 1 CI l3_2_0 [20] $end
$var wire 1 DI l3_2_0 [19] $end
$var wire 1 EI l3_2_0 [18] $end
$var wire 1 FI l3_2_0 [17] $end
$var wire 1 GI l3_2_0 [16] $end
$var wire 1 HI l3_2_0 [15] $end
$var wire 1 II l3_2_0 [14] $end
$var wire 1 JI l3_2_0 [13] $end
$var wire 1 KI l3_2_0 [12] $end
$var wire 1 LI l3_2_0 [11] $end
$var wire 1 MI l3_2_0 [10] $end
$var wire 1 NI l3_2_0 [9] $end
$var wire 1 OI l3_2_0 [8] $end
$var wire 1 PI l3_2_0 [7] $end
$var wire 1 QI l3_2_0 [6] $end
$var wire 1 RI l3_2_0 [5] $end
$var wire 1 SI l3_2_0 [4] $end
$var wire 1 TI l3_2_0 [3] $end
$var wire 1 UI l3_2_0 [2] $end
$var wire 1 VI l3_2_0 [1] $end
$var wire 1 WI l3_2_0 [0] $end
$var wire 1 XI l3_2_1 [54] $end
$var wire 1 YI l3_2_1 [53] $end
$var wire 1 ZI l3_2_1 [52] $end
$var wire 1 [I l3_2_1 [51] $end
$var wire 1 \I l3_2_1 [50] $end
$var wire 1 ]I l3_2_1 [49] $end
$var wire 1 ^I l3_2_1 [48] $end
$var wire 1 _I l3_2_1 [47] $end
$var wire 1 `I l3_2_1 [46] $end
$var wire 1 aI l3_2_1 [45] $end
$var wire 1 bI l3_2_1 [44] $end
$var wire 1 cI l3_2_1 [43] $end
$var wire 1 dI l3_2_1 [42] $end
$var wire 1 eI l3_2_1 [41] $end
$var wire 1 fI l3_2_1 [40] $end
$var wire 1 gI l3_2_1 [39] $end
$var wire 1 hI l3_2_1 [38] $end
$var wire 1 iI l3_2_1 [37] $end
$var wire 1 jI l3_2_1 [36] $end
$var wire 1 kI l3_2_1 [35] $end
$var wire 1 lI l3_2_1 [34] $end
$var wire 1 mI l3_2_1 [33] $end
$var wire 1 nI l3_2_1 [32] $end
$var wire 1 oI l3_2_1 [31] $end
$var wire 1 pI l3_2_1 [30] $end
$var wire 1 qI l3_2_1 [29] $end
$var wire 1 rI l3_2_1 [28] $end
$var wire 1 sI l3_2_1 [27] $end
$var wire 1 tI l3_2_1 [26] $end
$var wire 1 uI l3_2_1 [25] $end
$var wire 1 vI l3_2_1 [24] $end
$var wire 1 wI l3_2_1 [23] $end
$var wire 1 xI l3_2_1 [22] $end
$var wire 1 yI l3_2_1 [21] $end
$var wire 1 zI l3_2_1 [20] $end
$var wire 1 {I l3_2_1 [19] $end
$var wire 1 |I l3_2_1 [18] $end
$var wire 1 }I l3_2_1 [17] $end
$var wire 1 ~I l3_2_1 [16] $end
$var wire 1 !J l3_2_1 [15] $end
$var wire 1 "J l3_2_1 [14] $end
$var wire 1 #J l3_2_1 [13] $end
$var wire 1 $J l3_2_1 [12] $end
$var wire 1 %J l3_2_1 [11] $end
$var wire 1 &J l3_2_1 [10] $end
$var wire 1 'J l3_2_1 [9] $end
$var wire 1 (J l3_2_1 [8] $end
$var wire 1 )J l3_2_1 [7] $end
$var wire 1 *J l3_2_1 [6] $end
$var wire 1 +J l3_2_1 [5] $end
$var wire 1 ,J l3_2_1 [4] $end
$var wire 1 -J l3_2_1 [3] $end
$var wire 1 .J l3_2_1 [2] $end
$var wire 1 /J l3_2_1 [1] $end
$var wire 1 0J l3_2_1 [0] $end
$var wire 1 1J l3_2_2 [54] $end
$var wire 1 2J l3_2_2 [53] $end
$var wire 1 3J l3_2_2 [52] $end
$var wire 1 4J l3_2_2 [51] $end
$var wire 1 5J l3_2_2 [50] $end
$var wire 1 6J l3_2_2 [49] $end
$var wire 1 7J l3_2_2 [48] $end
$var wire 1 8J l3_2_2 [47] $end
$var wire 1 9J l3_2_2 [46] $end
$var wire 1 :J l3_2_2 [45] $end
$var wire 1 ;J l3_2_2 [44] $end
$var wire 1 <J l3_2_2 [43] $end
$var wire 1 =J l3_2_2 [42] $end
$var wire 1 >J l3_2_2 [41] $end
$var wire 1 ?J l3_2_2 [40] $end
$var wire 1 @J l3_2_2 [39] $end
$var wire 1 AJ l3_2_2 [38] $end
$var wire 1 BJ l3_2_2 [37] $end
$var wire 1 CJ l3_2_2 [36] $end
$var wire 1 DJ l3_2_2 [35] $end
$var wire 1 EJ l3_2_2 [34] $end
$var wire 1 FJ l3_2_2 [33] $end
$var wire 1 GJ l3_2_2 [32] $end
$var wire 1 HJ l3_2_2 [31] $end
$var wire 1 IJ l3_2_2 [30] $end
$var wire 1 JJ l3_2_2 [29] $end
$var wire 1 KJ l3_2_2 [28] $end
$var wire 1 LJ l3_2_2 [27] $end
$var wire 1 MJ l3_2_2 [26] $end
$var wire 1 NJ l3_2_2 [25] $end
$var wire 1 OJ l3_2_2 [24] $end
$var wire 1 PJ l3_2_2 [23] $end
$var wire 1 QJ l3_2_2 [22] $end
$var wire 1 RJ l3_2_2 [21] $end
$var wire 1 SJ l3_2_2 [20] $end
$var wire 1 TJ l3_2_2 [19] $end
$var wire 1 UJ l3_2_2 [18] $end
$var wire 1 VJ l3_2_2 [17] $end
$var wire 1 WJ l3_2_2 [16] $end
$var wire 1 XJ l3_2_2 [15] $end
$var wire 1 YJ l3_2_2 [14] $end
$var wire 1 ZJ l3_2_2 [13] $end
$var wire 1 [J l3_2_2 [12] $end
$var wire 1 \J l3_2_2 [11] $end
$var wire 1 ]J l3_2_2 [10] $end
$var wire 1 ^J l3_2_2 [9] $end
$var wire 1 _J l3_2_2 [8] $end
$var wire 1 `J l3_2_2 [7] $end
$var wire 1 aJ l3_2_2 [6] $end
$var wire 1 bJ l3_2_2 [5] $end
$var wire 1 cJ l3_2_2 [4] $end
$var wire 1 dJ l3_2_2 [3] $end
$var wire 1 eJ l3_2_2 [2] $end
$var wire 1 fJ l3_2_2 [1] $end
$var wire 1 gJ l3_2_2 [0] $end
$var wire 1 hJ l3_2_s [54] $end
$var wire 1 iJ l3_2_s [53] $end
$var wire 1 jJ l3_2_s [52] $end
$var wire 1 kJ l3_2_s [51] $end
$var wire 1 lJ l3_2_s [50] $end
$var wire 1 mJ l3_2_s [49] $end
$var wire 1 nJ l3_2_s [48] $end
$var wire 1 oJ l3_2_s [47] $end
$var wire 1 pJ l3_2_s [46] $end
$var wire 1 qJ l3_2_s [45] $end
$var wire 1 rJ l3_2_s [44] $end
$var wire 1 sJ l3_2_s [43] $end
$var wire 1 tJ l3_2_s [42] $end
$var wire 1 uJ l3_2_s [41] $end
$var wire 1 vJ l3_2_s [40] $end
$var wire 1 wJ l3_2_s [39] $end
$var wire 1 xJ l3_2_s [38] $end
$var wire 1 yJ l3_2_s [37] $end
$var wire 1 zJ l3_2_s [36] $end
$var wire 1 {J l3_2_s [35] $end
$var wire 1 |J l3_2_s [34] $end
$var wire 1 }J l3_2_s [33] $end
$var wire 1 ~J l3_2_s [32] $end
$var wire 1 !K l3_2_s [31] $end
$var wire 1 "K l3_2_s [30] $end
$var wire 1 #K l3_2_s [29] $end
$var wire 1 $K l3_2_s [28] $end
$var wire 1 %K l3_2_s [27] $end
$var wire 1 &K l3_2_s [26] $end
$var wire 1 'K l3_2_s [25] $end
$var wire 1 (K l3_2_s [24] $end
$var wire 1 )K l3_2_s [23] $end
$var wire 1 *K l3_2_s [22] $end
$var wire 1 +K l3_2_s [21] $end
$var wire 1 ,K l3_2_s [20] $end
$var wire 1 -K l3_2_s [19] $end
$var wire 1 .K l3_2_s [18] $end
$var wire 1 /K l3_2_s [17] $end
$var wire 1 0K l3_2_s [16] $end
$var wire 1 1K l3_2_s [15] $end
$var wire 1 2K l3_2_s [14] $end
$var wire 1 3K l3_2_s [13] $end
$var wire 1 4K l3_2_s [12] $end
$var wire 1 5K l3_2_s [11] $end
$var wire 1 6K l3_2_s [10] $end
$var wire 1 7K l3_2_s [9] $end
$var wire 1 8K l3_2_s [8] $end
$var wire 1 9K l3_2_s [7] $end
$var wire 1 :K l3_2_s [6] $end
$var wire 1 ;K l3_2_s [5] $end
$var wire 1 <K l3_2_s [4] $end
$var wire 1 =K l3_2_s [3] $end
$var wire 1 >K l3_2_s [2] $end
$var wire 1 ?K l3_2_s [1] $end
$var wire 1 @K l3_2_s [0] $end
$var wire 1 AK l3_2_ca [54] $end
$var wire 1 BK l3_2_ca [53] $end
$var wire 1 CK l3_2_ca [52] $end
$var wire 1 DK l3_2_ca [51] $end
$var wire 1 EK l3_2_ca [50] $end
$var wire 1 FK l3_2_ca [49] $end
$var wire 1 GK l3_2_ca [48] $end
$var wire 1 HK l3_2_ca [47] $end
$var wire 1 IK l3_2_ca [46] $end
$var wire 1 JK l3_2_ca [45] $end
$var wire 1 KK l3_2_ca [44] $end
$var wire 1 LK l3_2_ca [43] $end
$var wire 1 MK l3_2_ca [42] $end
$var wire 1 NK l3_2_ca [41] $end
$var wire 1 OK l3_2_ca [40] $end
$var wire 1 PK l3_2_ca [39] $end
$var wire 1 QK l3_2_ca [38] $end
$var wire 1 RK l3_2_ca [37] $end
$var wire 1 SK l3_2_ca [36] $end
$var wire 1 TK l3_2_ca [35] $end
$var wire 1 UK l3_2_ca [34] $end
$var wire 1 VK l3_2_ca [33] $end
$var wire 1 WK l3_2_ca [32] $end
$var wire 1 XK l3_2_ca [31] $end
$var wire 1 YK l3_2_ca [30] $end
$var wire 1 ZK l3_2_ca [29] $end
$var wire 1 [K l3_2_ca [28] $end
$var wire 1 \K l3_2_ca [27] $end
$var wire 1 ]K l3_2_ca [26] $end
$var wire 1 ^K l3_2_ca [25] $end
$var wire 1 _K l3_2_ca [24] $end
$var wire 1 `K l3_2_ca [23] $end
$var wire 1 aK l3_2_ca [22] $end
$var wire 1 bK l3_2_ca [21] $end
$var wire 1 cK l3_2_ca [20] $end
$var wire 1 dK l3_2_ca [19] $end
$var wire 1 eK l3_2_ca [18] $end
$var wire 1 fK l3_2_ca [17] $end
$var wire 1 gK l3_2_ca [16] $end
$var wire 1 hK l3_2_ca [15] $end
$var wire 1 iK l3_2_ca [14] $end
$var wire 1 jK l3_2_ca [13] $end
$var wire 1 kK l3_2_ca [12] $end
$var wire 1 lK l3_2_ca [11] $end
$var wire 1 mK l3_2_ca [10] $end
$var wire 1 nK l3_2_ca [9] $end
$var wire 1 oK l3_2_ca [8] $end
$var wire 1 pK l3_2_ca [7] $end
$var wire 1 qK l3_2_ca [6] $end
$var wire 1 rK l3_2_ca [5] $end
$var wire 1 sK l3_2_ca [4] $end
$var wire 1 tK l3_2_ca [3] $end
$var wire 1 uK l3_2_ca [2] $end
$var wire 1 vK l3_2_ca [1] $end
$var wire 1 wK l3_2_ca [0] $end
$var reg 55 xK l3_s1_reg [54:0] $end
$var reg 55 yK l3_c1_reg [54:0] $end
$var reg 55 zK l3_s2_reg [54:0] $end
$var reg 55 {K l3_c2_reg [54:0] $end
$var wire 1 |K l4_1_0 [63] $end
$var wire 1 }K l4_1_0 [62] $end
$var wire 1 ~K l4_1_0 [61] $end
$var wire 1 !L l4_1_0 [60] $end
$var wire 1 "L l4_1_0 [59] $end
$var wire 1 #L l4_1_0 [58] $end
$var wire 1 $L l4_1_0 [57] $end
$var wire 1 %L l4_1_0 [56] $end
$var wire 1 &L l4_1_0 [55] $end
$var wire 1 'L l4_1_0 [54] $end
$var wire 1 (L l4_1_0 [53] $end
$var wire 1 )L l4_1_0 [52] $end
$var wire 1 *L l4_1_0 [51] $end
$var wire 1 +L l4_1_0 [50] $end
$var wire 1 ,L l4_1_0 [49] $end
$var wire 1 -L l4_1_0 [48] $end
$var wire 1 .L l4_1_0 [47] $end
$var wire 1 /L l4_1_0 [46] $end
$var wire 1 0L l4_1_0 [45] $end
$var wire 1 1L l4_1_0 [44] $end
$var wire 1 2L l4_1_0 [43] $end
$var wire 1 3L l4_1_0 [42] $end
$var wire 1 4L l4_1_0 [41] $end
$var wire 1 5L l4_1_0 [40] $end
$var wire 1 6L l4_1_0 [39] $end
$var wire 1 7L l4_1_0 [38] $end
$var wire 1 8L l4_1_0 [37] $end
$var wire 1 9L l4_1_0 [36] $end
$var wire 1 :L l4_1_0 [35] $end
$var wire 1 ;L l4_1_0 [34] $end
$var wire 1 <L l4_1_0 [33] $end
$var wire 1 =L l4_1_0 [32] $end
$var wire 1 >L l4_1_0 [31] $end
$var wire 1 ?L l4_1_0 [30] $end
$var wire 1 @L l4_1_0 [29] $end
$var wire 1 AL l4_1_0 [28] $end
$var wire 1 BL l4_1_0 [27] $end
$var wire 1 CL l4_1_0 [26] $end
$var wire 1 DL l4_1_0 [25] $end
$var wire 1 EL l4_1_0 [24] $end
$var wire 1 FL l4_1_0 [23] $end
$var wire 1 GL l4_1_0 [22] $end
$var wire 1 HL l4_1_0 [21] $end
$var wire 1 IL l4_1_0 [20] $end
$var wire 1 JL l4_1_0 [19] $end
$var wire 1 KL l4_1_0 [18] $end
$var wire 1 LL l4_1_0 [17] $end
$var wire 1 ML l4_1_0 [16] $end
$var wire 1 NL l4_1_0 [15] $end
$var wire 1 OL l4_1_0 [14] $end
$var wire 1 PL l4_1_0 [13] $end
$var wire 1 QL l4_1_0 [12] $end
$var wire 1 RL l4_1_0 [11] $end
$var wire 1 SL l4_1_0 [10] $end
$var wire 1 TL l4_1_0 [9] $end
$var wire 1 UL l4_1_0 [8] $end
$var wire 1 VL l4_1_0 [7] $end
$var wire 1 WL l4_1_0 [6] $end
$var wire 1 XL l4_1_0 [5] $end
$var wire 1 YL l4_1_0 [4] $end
$var wire 1 ZL l4_1_0 [3] $end
$var wire 1 [L l4_1_0 [2] $end
$var wire 1 \L l4_1_0 [1] $end
$var wire 1 ]L l4_1_0 [0] $end
$var wire 1 ^L l4_1_1 [63] $end
$var wire 1 _L l4_1_1 [62] $end
$var wire 1 `L l4_1_1 [61] $end
$var wire 1 aL l4_1_1 [60] $end
$var wire 1 bL l4_1_1 [59] $end
$var wire 1 cL l4_1_1 [58] $end
$var wire 1 dL l4_1_1 [57] $end
$var wire 1 eL l4_1_1 [56] $end
$var wire 1 fL l4_1_1 [55] $end
$var wire 1 gL l4_1_1 [54] $end
$var wire 1 hL l4_1_1 [53] $end
$var wire 1 iL l4_1_1 [52] $end
$var wire 1 jL l4_1_1 [51] $end
$var wire 1 kL l4_1_1 [50] $end
$var wire 1 lL l4_1_1 [49] $end
$var wire 1 mL l4_1_1 [48] $end
$var wire 1 nL l4_1_1 [47] $end
$var wire 1 oL l4_1_1 [46] $end
$var wire 1 pL l4_1_1 [45] $end
$var wire 1 qL l4_1_1 [44] $end
$var wire 1 rL l4_1_1 [43] $end
$var wire 1 sL l4_1_1 [42] $end
$var wire 1 tL l4_1_1 [41] $end
$var wire 1 uL l4_1_1 [40] $end
$var wire 1 vL l4_1_1 [39] $end
$var wire 1 wL l4_1_1 [38] $end
$var wire 1 xL l4_1_1 [37] $end
$var wire 1 yL l4_1_1 [36] $end
$var wire 1 zL l4_1_1 [35] $end
$var wire 1 {L l4_1_1 [34] $end
$var wire 1 |L l4_1_1 [33] $end
$var wire 1 }L l4_1_1 [32] $end
$var wire 1 ~L l4_1_1 [31] $end
$var wire 1 !M l4_1_1 [30] $end
$var wire 1 "M l4_1_1 [29] $end
$var wire 1 #M l4_1_1 [28] $end
$var wire 1 $M l4_1_1 [27] $end
$var wire 1 %M l4_1_1 [26] $end
$var wire 1 &M l4_1_1 [25] $end
$var wire 1 'M l4_1_1 [24] $end
$var wire 1 (M l4_1_1 [23] $end
$var wire 1 )M l4_1_1 [22] $end
$var wire 1 *M l4_1_1 [21] $end
$var wire 1 +M l4_1_1 [20] $end
$var wire 1 ,M l4_1_1 [19] $end
$var wire 1 -M l4_1_1 [18] $end
$var wire 1 .M l4_1_1 [17] $end
$var wire 1 /M l4_1_1 [16] $end
$var wire 1 0M l4_1_1 [15] $end
$var wire 1 1M l4_1_1 [14] $end
$var wire 1 2M l4_1_1 [13] $end
$var wire 1 3M l4_1_1 [12] $end
$var wire 1 4M l4_1_1 [11] $end
$var wire 1 5M l4_1_1 [10] $end
$var wire 1 6M l4_1_1 [9] $end
$var wire 1 7M l4_1_1 [8] $end
$var wire 1 8M l4_1_1 [7] $end
$var wire 1 9M l4_1_1 [6] $end
$var wire 1 :M l4_1_1 [5] $end
$var wire 1 ;M l4_1_1 [4] $end
$var wire 1 <M l4_1_1 [3] $end
$var wire 1 =M l4_1_1 [2] $end
$var wire 1 >M l4_1_1 [1] $end
$var wire 1 ?M l4_1_1 [0] $end
$var wire 1 @M l4_1_2 [63] $end
$var wire 1 AM l4_1_2 [62] $end
$var wire 1 BM l4_1_2 [61] $end
$var wire 1 CM l4_1_2 [60] $end
$var wire 1 DM l4_1_2 [59] $end
$var wire 1 EM l4_1_2 [58] $end
$var wire 1 FM l4_1_2 [57] $end
$var wire 1 GM l4_1_2 [56] $end
$var wire 1 HM l4_1_2 [55] $end
$var wire 1 IM l4_1_2 [54] $end
$var wire 1 JM l4_1_2 [53] $end
$var wire 1 KM l4_1_2 [52] $end
$var wire 1 LM l4_1_2 [51] $end
$var wire 1 MM l4_1_2 [50] $end
$var wire 1 NM l4_1_2 [49] $end
$var wire 1 OM l4_1_2 [48] $end
$var wire 1 PM l4_1_2 [47] $end
$var wire 1 QM l4_1_2 [46] $end
$var wire 1 RM l4_1_2 [45] $end
$var wire 1 SM l4_1_2 [44] $end
$var wire 1 TM l4_1_2 [43] $end
$var wire 1 UM l4_1_2 [42] $end
$var wire 1 VM l4_1_2 [41] $end
$var wire 1 WM l4_1_2 [40] $end
$var wire 1 XM l4_1_2 [39] $end
$var wire 1 YM l4_1_2 [38] $end
$var wire 1 ZM l4_1_2 [37] $end
$var wire 1 [M l4_1_2 [36] $end
$var wire 1 \M l4_1_2 [35] $end
$var wire 1 ]M l4_1_2 [34] $end
$var wire 1 ^M l4_1_2 [33] $end
$var wire 1 _M l4_1_2 [32] $end
$var wire 1 `M l4_1_2 [31] $end
$var wire 1 aM l4_1_2 [30] $end
$var wire 1 bM l4_1_2 [29] $end
$var wire 1 cM l4_1_2 [28] $end
$var wire 1 dM l4_1_2 [27] $end
$var wire 1 eM l4_1_2 [26] $end
$var wire 1 fM l4_1_2 [25] $end
$var wire 1 gM l4_1_2 [24] $end
$var wire 1 hM l4_1_2 [23] $end
$var wire 1 iM l4_1_2 [22] $end
$var wire 1 jM l4_1_2 [21] $end
$var wire 1 kM l4_1_2 [20] $end
$var wire 1 lM l4_1_2 [19] $end
$var wire 1 mM l4_1_2 [18] $end
$var wire 1 nM l4_1_2 [17] $end
$var wire 1 oM l4_1_2 [16] $end
$var wire 1 pM l4_1_2 [15] $end
$var wire 1 qM l4_1_2 [14] $end
$var wire 1 rM l4_1_2 [13] $end
$var wire 1 sM l4_1_2 [12] $end
$var wire 1 tM l4_1_2 [11] $end
$var wire 1 uM l4_1_2 [10] $end
$var wire 1 vM l4_1_2 [9] $end
$var wire 1 wM l4_1_2 [8] $end
$var wire 1 xM l4_1_2 [7] $end
$var wire 1 yM l4_1_2 [6] $end
$var wire 1 zM l4_1_2 [5] $end
$var wire 1 {M l4_1_2 [4] $end
$var wire 1 |M l4_1_2 [3] $end
$var wire 1 }M l4_1_2 [2] $end
$var wire 1 ~M l4_1_2 [1] $end
$var wire 1 !N l4_1_2 [0] $end
$var wire 1 "N l4_1_3 [63] $end
$var wire 1 #N l4_1_3 [62] $end
$var wire 1 $N l4_1_3 [61] $end
$var wire 1 %N l4_1_3 [60] $end
$var wire 1 &N l4_1_3 [59] $end
$var wire 1 'N l4_1_3 [58] $end
$var wire 1 (N l4_1_3 [57] $end
$var wire 1 )N l4_1_3 [56] $end
$var wire 1 *N l4_1_3 [55] $end
$var wire 1 +N l4_1_3 [54] $end
$var wire 1 ,N l4_1_3 [53] $end
$var wire 1 -N l4_1_3 [52] $end
$var wire 1 .N l4_1_3 [51] $end
$var wire 1 /N l4_1_3 [50] $end
$var wire 1 0N l4_1_3 [49] $end
$var wire 1 1N l4_1_3 [48] $end
$var wire 1 2N l4_1_3 [47] $end
$var wire 1 3N l4_1_3 [46] $end
$var wire 1 4N l4_1_3 [45] $end
$var wire 1 5N l4_1_3 [44] $end
$var wire 1 6N l4_1_3 [43] $end
$var wire 1 7N l4_1_3 [42] $end
$var wire 1 8N l4_1_3 [41] $end
$var wire 1 9N l4_1_3 [40] $end
$var wire 1 :N l4_1_3 [39] $end
$var wire 1 ;N l4_1_3 [38] $end
$var wire 1 <N l4_1_3 [37] $end
$var wire 1 =N l4_1_3 [36] $end
$var wire 1 >N l4_1_3 [35] $end
$var wire 1 ?N l4_1_3 [34] $end
$var wire 1 @N l4_1_3 [33] $end
$var wire 1 AN l4_1_3 [32] $end
$var wire 1 BN l4_1_3 [31] $end
$var wire 1 CN l4_1_3 [30] $end
$var wire 1 DN l4_1_3 [29] $end
$var wire 1 EN l4_1_3 [28] $end
$var wire 1 FN l4_1_3 [27] $end
$var wire 1 GN l4_1_3 [26] $end
$var wire 1 HN l4_1_3 [25] $end
$var wire 1 IN l4_1_3 [24] $end
$var wire 1 JN l4_1_3 [23] $end
$var wire 1 KN l4_1_3 [22] $end
$var wire 1 LN l4_1_3 [21] $end
$var wire 1 MN l4_1_3 [20] $end
$var wire 1 NN l4_1_3 [19] $end
$var wire 1 ON l4_1_3 [18] $end
$var wire 1 PN l4_1_3 [17] $end
$var wire 1 QN l4_1_3 [16] $end
$var wire 1 RN l4_1_3 [15] $end
$var wire 1 SN l4_1_3 [14] $end
$var wire 1 TN l4_1_3 [13] $end
$var wire 1 UN l4_1_3 [12] $end
$var wire 1 VN l4_1_3 [11] $end
$var wire 1 WN l4_1_3 [10] $end
$var wire 1 XN l4_1_3 [9] $end
$var wire 1 YN l4_1_3 [8] $end
$var wire 1 ZN l4_1_3 [7] $end
$var wire 1 [N l4_1_3 [6] $end
$var wire 1 \N l4_1_3 [5] $end
$var wire 1 ]N l4_1_3 [4] $end
$var wire 1 ^N l4_1_3 [3] $end
$var wire 1 _N l4_1_3 [2] $end
$var wire 1 `N l4_1_3 [1] $end
$var wire 1 aN l4_1_3 [0] $end
$var wire 1 bN l4_1_s [63] $end
$var wire 1 cN l4_1_s [62] $end
$var wire 1 dN l4_1_s [61] $end
$var wire 1 eN l4_1_s [60] $end
$var wire 1 fN l4_1_s [59] $end
$var wire 1 gN l4_1_s [58] $end
$var wire 1 hN l4_1_s [57] $end
$var wire 1 iN l4_1_s [56] $end
$var wire 1 jN l4_1_s [55] $end
$var wire 1 kN l4_1_s [54] $end
$var wire 1 lN l4_1_s [53] $end
$var wire 1 mN l4_1_s [52] $end
$var wire 1 nN l4_1_s [51] $end
$var wire 1 oN l4_1_s [50] $end
$var wire 1 pN l4_1_s [49] $end
$var wire 1 qN l4_1_s [48] $end
$var wire 1 rN l4_1_s [47] $end
$var wire 1 sN l4_1_s [46] $end
$var wire 1 tN l4_1_s [45] $end
$var wire 1 uN l4_1_s [44] $end
$var wire 1 vN l4_1_s [43] $end
$var wire 1 wN l4_1_s [42] $end
$var wire 1 xN l4_1_s [41] $end
$var wire 1 yN l4_1_s [40] $end
$var wire 1 zN l4_1_s [39] $end
$var wire 1 {N l4_1_s [38] $end
$var wire 1 |N l4_1_s [37] $end
$var wire 1 }N l4_1_s [36] $end
$var wire 1 ~N l4_1_s [35] $end
$var wire 1 !O l4_1_s [34] $end
$var wire 1 "O l4_1_s [33] $end
$var wire 1 #O l4_1_s [32] $end
$var wire 1 $O l4_1_s [31] $end
$var wire 1 %O l4_1_s [30] $end
$var wire 1 &O l4_1_s [29] $end
$var wire 1 'O l4_1_s [28] $end
$var wire 1 (O l4_1_s [27] $end
$var wire 1 )O l4_1_s [26] $end
$var wire 1 *O l4_1_s [25] $end
$var wire 1 +O l4_1_s [24] $end
$var wire 1 ,O l4_1_s [23] $end
$var wire 1 -O l4_1_s [22] $end
$var wire 1 .O l4_1_s [21] $end
$var wire 1 /O l4_1_s [20] $end
$var wire 1 0O l4_1_s [19] $end
$var wire 1 1O l4_1_s [18] $end
$var wire 1 2O l4_1_s [17] $end
$var wire 1 3O l4_1_s [16] $end
$var wire 1 4O l4_1_s [15] $end
$var wire 1 5O l4_1_s [14] $end
$var wire 1 6O l4_1_s [13] $end
$var wire 1 7O l4_1_s [12] $end
$var wire 1 8O l4_1_s [11] $end
$var wire 1 9O l4_1_s [10] $end
$var wire 1 :O l4_1_s [9] $end
$var wire 1 ;O l4_1_s [8] $end
$var wire 1 <O l4_1_s [7] $end
$var wire 1 =O l4_1_s [6] $end
$var wire 1 >O l4_1_s [5] $end
$var wire 1 ?O l4_1_s [4] $end
$var wire 1 @O l4_1_s [3] $end
$var wire 1 AO l4_1_s [2] $end
$var wire 1 BO l4_1_s [1] $end
$var wire 1 CO l4_1_s [0] $end
$var wire 1 DO l4_1_ca [63] $end
$var wire 1 EO l4_1_ca [62] $end
$var wire 1 FO l4_1_ca [61] $end
$var wire 1 GO l4_1_ca [60] $end
$var wire 1 HO l4_1_ca [59] $end
$var wire 1 IO l4_1_ca [58] $end
$var wire 1 JO l4_1_ca [57] $end
$var wire 1 KO l4_1_ca [56] $end
$var wire 1 LO l4_1_ca [55] $end
$var wire 1 MO l4_1_ca [54] $end
$var wire 1 NO l4_1_ca [53] $end
$var wire 1 OO l4_1_ca [52] $end
$var wire 1 PO l4_1_ca [51] $end
$var wire 1 QO l4_1_ca [50] $end
$var wire 1 RO l4_1_ca [49] $end
$var wire 1 SO l4_1_ca [48] $end
$var wire 1 TO l4_1_ca [47] $end
$var wire 1 UO l4_1_ca [46] $end
$var wire 1 VO l4_1_ca [45] $end
$var wire 1 WO l4_1_ca [44] $end
$var wire 1 XO l4_1_ca [43] $end
$var wire 1 YO l4_1_ca [42] $end
$var wire 1 ZO l4_1_ca [41] $end
$var wire 1 [O l4_1_ca [40] $end
$var wire 1 \O l4_1_ca [39] $end
$var wire 1 ]O l4_1_ca [38] $end
$var wire 1 ^O l4_1_ca [37] $end
$var wire 1 _O l4_1_ca [36] $end
$var wire 1 `O l4_1_ca [35] $end
$var wire 1 aO l4_1_ca [34] $end
$var wire 1 bO l4_1_ca [33] $end
$var wire 1 cO l4_1_ca [32] $end
$var wire 1 dO l4_1_ca [31] $end
$var wire 1 eO l4_1_ca [30] $end
$var wire 1 fO l4_1_ca [29] $end
$var wire 1 gO l4_1_ca [28] $end
$var wire 1 hO l4_1_ca [27] $end
$var wire 1 iO l4_1_ca [26] $end
$var wire 1 jO l4_1_ca [25] $end
$var wire 1 kO l4_1_ca [24] $end
$var wire 1 lO l4_1_ca [23] $end
$var wire 1 mO l4_1_ca [22] $end
$var wire 1 nO l4_1_ca [21] $end
$var wire 1 oO l4_1_ca [20] $end
$var wire 1 pO l4_1_ca [19] $end
$var wire 1 qO l4_1_ca [18] $end
$var wire 1 rO l4_1_ca [17] $end
$var wire 1 sO l4_1_ca [16] $end
$var wire 1 tO l4_1_ca [15] $end
$var wire 1 uO l4_1_ca [14] $end
$var wire 1 vO l4_1_ca [13] $end
$var wire 1 wO l4_1_ca [12] $end
$var wire 1 xO l4_1_ca [11] $end
$var wire 1 yO l4_1_ca [10] $end
$var wire 1 zO l4_1_ca [9] $end
$var wire 1 {O l4_1_ca [8] $end
$var wire 1 |O l4_1_ca [7] $end
$var wire 1 }O l4_1_ca [6] $end
$var wire 1 ~O l4_1_ca [5] $end
$var wire 1 !P l4_1_ca [4] $end
$var wire 1 "P l4_1_ca [3] $end
$var wire 1 #P l4_1_ca [2] $end
$var wire 1 $P l4_1_ca [1] $end
$var wire 1 %P l4_1_ca [0] $end
$var wire 1 &P l4_1_cin [63] $end
$var wire 1 'P l4_1_cin [62] $end
$var wire 1 (P l4_1_cin [61] $end
$var wire 1 )P l4_1_cin [60] $end
$var wire 1 *P l4_1_cin [59] $end
$var wire 1 +P l4_1_cin [58] $end
$var wire 1 ,P l4_1_cin [57] $end
$var wire 1 -P l4_1_cin [56] $end
$var wire 1 .P l4_1_cin [55] $end
$var wire 1 /P l4_1_cin [54] $end
$var wire 1 0P l4_1_cin [53] $end
$var wire 1 1P l4_1_cin [52] $end
$var wire 1 2P l4_1_cin [51] $end
$var wire 1 3P l4_1_cin [50] $end
$var wire 1 4P l4_1_cin [49] $end
$var wire 1 5P l4_1_cin [48] $end
$var wire 1 6P l4_1_cin [47] $end
$var wire 1 7P l4_1_cin [46] $end
$var wire 1 8P l4_1_cin [45] $end
$var wire 1 9P l4_1_cin [44] $end
$var wire 1 :P l4_1_cin [43] $end
$var wire 1 ;P l4_1_cin [42] $end
$var wire 1 <P l4_1_cin [41] $end
$var wire 1 =P l4_1_cin [40] $end
$var wire 1 >P l4_1_cin [39] $end
$var wire 1 ?P l4_1_cin [38] $end
$var wire 1 @P l4_1_cin [37] $end
$var wire 1 AP l4_1_cin [36] $end
$var wire 1 BP l4_1_cin [35] $end
$var wire 1 CP l4_1_cin [34] $end
$var wire 1 DP l4_1_cin [33] $end
$var wire 1 EP l4_1_cin [32] $end
$var wire 1 FP l4_1_cin [31] $end
$var wire 1 GP l4_1_cin [30] $end
$var wire 1 HP l4_1_cin [29] $end
$var wire 1 IP l4_1_cin [28] $end
$var wire 1 JP l4_1_cin [27] $end
$var wire 1 KP l4_1_cin [26] $end
$var wire 1 LP l4_1_cin [25] $end
$var wire 1 MP l4_1_cin [24] $end
$var wire 1 NP l4_1_cin [23] $end
$var wire 1 OP l4_1_cin [22] $end
$var wire 1 PP l4_1_cin [21] $end
$var wire 1 QP l4_1_cin [20] $end
$var wire 1 RP l4_1_cin [19] $end
$var wire 1 SP l4_1_cin [18] $end
$var wire 1 TP l4_1_cin [17] $end
$var wire 1 UP l4_1_cin [16] $end
$var wire 1 VP l4_1_cin [15] $end
$var wire 1 WP l4_1_cin [14] $end
$var wire 1 XP l4_1_cin [13] $end
$var wire 1 YP l4_1_cin [12] $end
$var wire 1 ZP l4_1_cin [11] $end
$var wire 1 [P l4_1_cin [10] $end
$var wire 1 \P l4_1_cin [9] $end
$var wire 1 ]P l4_1_cin [8] $end
$var wire 1 ^P l4_1_cin [7] $end
$var wire 1 _P l4_1_cin [6] $end
$var wire 1 `P l4_1_cin [5] $end
$var wire 1 aP l4_1_cin [4] $end
$var wire 1 bP l4_1_cin [3] $end
$var wire 1 cP l4_1_cin [2] $end
$var wire 1 dP l4_1_cin [1] $end
$var wire 1 eP l4_1_cin [0] $end
$var wire 1 fP l4_1_cout [63] $end
$var wire 1 gP l4_1_cout [62] $end
$var wire 1 hP l4_1_cout [61] $end
$var wire 1 iP l4_1_cout [60] $end
$var wire 1 jP l4_1_cout [59] $end
$var wire 1 kP l4_1_cout [58] $end
$var wire 1 lP l4_1_cout [57] $end
$var wire 1 mP l4_1_cout [56] $end
$var wire 1 nP l4_1_cout [55] $end
$var wire 1 oP l4_1_cout [54] $end
$var wire 1 pP l4_1_cout [53] $end
$var wire 1 qP l4_1_cout [52] $end
$var wire 1 rP l4_1_cout [51] $end
$var wire 1 sP l4_1_cout [50] $end
$var wire 1 tP l4_1_cout [49] $end
$var wire 1 uP l4_1_cout [48] $end
$var wire 1 vP l4_1_cout [47] $end
$var wire 1 wP l4_1_cout [46] $end
$var wire 1 xP l4_1_cout [45] $end
$var wire 1 yP l4_1_cout [44] $end
$var wire 1 zP l4_1_cout [43] $end
$var wire 1 {P l4_1_cout [42] $end
$var wire 1 |P l4_1_cout [41] $end
$var wire 1 }P l4_1_cout [40] $end
$var wire 1 ~P l4_1_cout [39] $end
$var wire 1 !Q l4_1_cout [38] $end
$var wire 1 "Q l4_1_cout [37] $end
$var wire 1 #Q l4_1_cout [36] $end
$var wire 1 $Q l4_1_cout [35] $end
$var wire 1 %Q l4_1_cout [34] $end
$var wire 1 &Q l4_1_cout [33] $end
$var wire 1 'Q l4_1_cout [32] $end
$var wire 1 (Q l4_1_cout [31] $end
$var wire 1 )Q l4_1_cout [30] $end
$var wire 1 *Q l4_1_cout [29] $end
$var wire 1 +Q l4_1_cout [28] $end
$var wire 1 ,Q l4_1_cout [27] $end
$var wire 1 -Q l4_1_cout [26] $end
$var wire 1 .Q l4_1_cout [25] $end
$var wire 1 /Q l4_1_cout [24] $end
$var wire 1 0Q l4_1_cout [23] $end
$var wire 1 1Q l4_1_cout [22] $end
$var wire 1 2Q l4_1_cout [21] $end
$var wire 1 3Q l4_1_cout [20] $end
$var wire 1 4Q l4_1_cout [19] $end
$var wire 1 5Q l4_1_cout [18] $end
$var wire 1 6Q l4_1_cout [17] $end
$var wire 1 7Q l4_1_cout [16] $end
$var wire 1 8Q l4_1_cout [15] $end
$var wire 1 9Q l4_1_cout [14] $end
$var wire 1 :Q l4_1_cout [13] $end
$var wire 1 ;Q l4_1_cout [12] $end
$var wire 1 <Q l4_1_cout [11] $end
$var wire 1 =Q l4_1_cout [10] $end
$var wire 1 >Q l4_1_cout [9] $end
$var wire 1 ?Q l4_1_cout [8] $end
$var wire 1 @Q l4_1_cout [7] $end
$var wire 1 AQ l4_1_cout [6] $end
$var wire 1 BQ l4_1_cout [5] $end
$var wire 1 CQ l4_1_cout [4] $end
$var wire 1 DQ l4_1_cout [3] $end
$var wire 1 EQ l4_1_cout [2] $end
$var wire 1 FQ l4_1_cout [1] $end
$var wire 1 GQ l4_1_cout [0] $end
$var reg 64 HQ s [63:0] $end
$var reg 64 IQ c [63:0] $end

$scope module boothcode0 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 6" code [2] $end
$var wire 1 7" code [1] $end
$var wire 1 JQ code [0] $end
$var reg 33 KQ product [32:0] $end
$var reg 2 LQ h [1:0] $end
$var reg 1 MQ s $end
$upscope $end

$scope module boothcode1 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 4" code [2] $end
$var wire 1 5" code [1] $end
$var wire 1 6" code [0] $end
$var reg 33 NQ product [32:0] $end
$var reg 2 OQ h [1:0] $end
$var reg 1 PQ s $end
$upscope $end

$scope module boothcode2 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 2" code [2] $end
$var wire 1 3" code [1] $end
$var wire 1 4" code [0] $end
$var reg 33 QQ product [32:0] $end
$var reg 2 RQ h [1:0] $end
$var reg 1 SQ s $end
$upscope $end

$scope module boothcode3 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 0" code [2] $end
$var wire 1 1" code [1] $end
$var wire 1 2" code [0] $end
$var reg 33 TQ product [32:0] $end
$var reg 2 UQ h [1:0] $end
$var reg 1 VQ s $end
$upscope $end

$scope module boothcode4 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 ." code [2] $end
$var wire 1 /" code [1] $end
$var wire 1 0" code [0] $end
$var reg 33 WQ product [32:0] $end
$var reg 2 XQ h [1:0] $end
$var reg 1 YQ s $end
$upscope $end

$scope module boothcode5 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 ," code [2] $end
$var wire 1 -" code [1] $end
$var wire 1 ." code [0] $end
$var reg 33 ZQ product [32:0] $end
$var reg 2 [Q h [1:0] $end
$var reg 1 \Q s $end
$upscope $end

$scope module boothcode6 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 *" code [2] $end
$var wire 1 +" code [1] $end
$var wire 1 ," code [0] $end
$var reg 33 ]Q product [32:0] $end
$var reg 2 ^Q h [1:0] $end
$var reg 1 _Q s $end
$upscope $end

$scope module boothcode7 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 (" code [2] $end
$var wire 1 )" code [1] $end
$var wire 1 *" code [0] $end
$var reg 33 `Q product [32:0] $end
$var reg 2 aQ h [1:0] $end
$var reg 1 bQ s $end
$upscope $end

$scope module boothcode8 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 &" code [2] $end
$var wire 1 '" code [1] $end
$var wire 1 (" code [0] $end
$var reg 33 cQ product [32:0] $end
$var reg 2 dQ h [1:0] $end
$var reg 1 eQ s $end
$upscope $end

$scope module boothcode9 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 $" code [2] $end
$var wire 1 %" code [1] $end
$var wire 1 &" code [0] $end
$var reg 33 fQ product [32:0] $end
$var reg 2 gQ h [1:0] $end
$var reg 1 hQ s $end
$upscope $end

$scope module boothcode10 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 "" code [2] $end
$var wire 1 #" code [1] $end
$var wire 1 $" code [0] $end
$var reg 33 iQ product [32:0] $end
$var reg 2 jQ h [1:0] $end
$var reg 1 kQ s $end
$upscope $end

$scope module boothcode11 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 ~! code [2] $end
$var wire 1 !" code [1] $end
$var wire 1 "" code [0] $end
$var reg 33 lQ product [32:0] $end
$var reg 2 mQ h [1:0] $end
$var reg 1 nQ s $end
$upscope $end

$scope module boothcode12 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 |! code [2] $end
$var wire 1 }! code [1] $end
$var wire 1 ~! code [0] $end
$var reg 33 oQ product [32:0] $end
$var reg 2 pQ h [1:0] $end
$var reg 1 qQ s $end
$upscope $end

$scope module boothcode13 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 z! code [2] $end
$var wire 1 {! code [1] $end
$var wire 1 |! code [0] $end
$var reg 33 rQ product [32:0] $end
$var reg 2 sQ h [1:0] $end
$var reg 1 tQ s $end
$upscope $end

$scope module boothcode14 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 x! code [2] $end
$var wire 1 y! code [1] $end
$var wire 1 z! code [0] $end
$var reg 33 uQ product [32:0] $end
$var reg 2 vQ h [1:0] $end
$var reg 1 wQ s $end
$upscope $end

$scope module boothcode15 $end
$var wire 1 S( A [31] $end
$var wire 1 T( A [30] $end
$var wire 1 U( A [29] $end
$var wire 1 V( A [28] $end
$var wire 1 W( A [27] $end
$var wire 1 X( A [26] $end
$var wire 1 Y( A [25] $end
$var wire 1 Z( A [24] $end
$var wire 1 [( A [23] $end
$var wire 1 \( A [22] $end
$var wire 1 ]( A [21] $end
$var wire 1 ^( A [20] $end
$var wire 1 _( A [19] $end
$var wire 1 `( A [18] $end
$var wire 1 a( A [17] $end
$var wire 1 b( A [16] $end
$var wire 1 c( A [15] $end
$var wire 1 d( A [14] $end
$var wire 1 e( A [13] $end
$var wire 1 f( A [12] $end
$var wire 1 g( A [11] $end
$var wire 1 h( A [10] $end
$var wire 1 i( A [9] $end
$var wire 1 j( A [8] $end
$var wire 1 k( A [7] $end
$var wire 1 l( A [6] $end
$var wire 1 m( A [5] $end
$var wire 1 n( A [4] $end
$var wire 1 o( A [3] $end
$var wire 1 p( A [2] $end
$var wire 1 q( A [1] $end
$var wire 1 r( A [0] $end
$var wire 1 v! code [2] $end
$var wire 1 w! code [1] $end
$var wire 1 x! code [0] $end
$var reg 33 xQ product [32:0] $end
$var reg 2 yQ h [1:0] $end
$var reg 1 zQ s $end
$upscope $end

$scope module l1_1 $end
$var parameter 32 {Q size $end
$var wire 1 &) c0 [35] $end
$var wire 1 ') c0 [34] $end
$var wire 1 () c0 [33] $end
$var wire 1 )) c0 [32] $end
$var wire 1 *) c0 [31] $end
$var wire 1 +) c0 [30] $end
$var wire 1 ,) c0 [29] $end
$var wire 1 -) c0 [28] $end
$var wire 1 .) c0 [27] $end
$var wire 1 /) c0 [26] $end
$var wire 1 0) c0 [25] $end
$var wire 1 1) c0 [24] $end
$var wire 1 2) c0 [23] $end
$var wire 1 3) c0 [22] $end
$var wire 1 4) c0 [21] $end
$var wire 1 5) c0 [20] $end
$var wire 1 6) c0 [19] $end
$var wire 1 7) c0 [18] $end
$var wire 1 8) c0 [17] $end
$var wire 1 9) c0 [16] $end
$var wire 1 :) c0 [15] $end
$var wire 1 ;) c0 [14] $end
$var wire 1 <) c0 [13] $end
$var wire 1 =) c0 [12] $end
$var wire 1 >) c0 [11] $end
$var wire 1 ?) c0 [10] $end
$var wire 1 @) c0 [9] $end
$var wire 1 A) c0 [8] $end
$var wire 1 B) c0 [7] $end
$var wire 1 C) c0 [6] $end
$var wire 1 D) c0 [5] $end
$var wire 1 E) c0 [4] $end
$var wire 1 F) c0 [3] $end
$var wire 1 G) c0 [2] $end
$var wire 1 H) c0 [1] $end
$var wire 1 I) c0 [0] $end
$var wire 1 J) c1 [35] $end
$var wire 1 K) c1 [34] $end
$var wire 1 L) c1 [33] $end
$var wire 1 M) c1 [32] $end
$var wire 1 N) c1 [31] $end
$var wire 1 O) c1 [30] $end
$var wire 1 P) c1 [29] $end
$var wire 1 Q) c1 [28] $end
$var wire 1 R) c1 [27] $end
$var wire 1 S) c1 [26] $end
$var wire 1 T) c1 [25] $end
$var wire 1 U) c1 [24] $end
$var wire 1 V) c1 [23] $end
$var wire 1 W) c1 [22] $end
$var wire 1 X) c1 [21] $end
$var wire 1 Y) c1 [20] $end
$var wire 1 Z) c1 [19] $end
$var wire 1 [) c1 [18] $end
$var wire 1 \) c1 [17] $end
$var wire 1 ]) c1 [16] $end
$var wire 1 ^) c1 [15] $end
$var wire 1 _) c1 [14] $end
$var wire 1 `) c1 [13] $end
$var wire 1 a) c1 [12] $end
$var wire 1 b) c1 [11] $end
$var wire 1 c) c1 [10] $end
$var wire 1 d) c1 [9] $end
$var wire 1 e) c1 [8] $end
$var wire 1 f) c1 [7] $end
$var wire 1 g) c1 [6] $end
$var wire 1 h) c1 [5] $end
$var wire 1 i) c1 [4] $end
$var wire 1 j) c1 [3] $end
$var wire 1 k) c1 [2] $end
$var wire 1 l) c1 [1] $end
$var wire 1 m) c1 [0] $end
$var wire 1 n) c2 [35] $end
$var wire 1 o) c2 [34] $end
$var wire 1 p) c2 [33] $end
$var wire 1 q) c2 [32] $end
$var wire 1 r) c2 [31] $end
$var wire 1 s) c2 [30] $end
$var wire 1 t) c2 [29] $end
$var wire 1 u) c2 [28] $end
$var wire 1 v) c2 [27] $end
$var wire 1 w) c2 [26] $end
$var wire 1 x) c2 [25] $end
$var wire 1 y) c2 [24] $end
$var wire 1 z) c2 [23] $end
$var wire 1 {) c2 [22] $end
$var wire 1 |) c2 [21] $end
$var wire 1 }) c2 [20] $end
$var wire 1 ~) c2 [19] $end
$var wire 1 !* c2 [18] $end
$var wire 1 "* c2 [17] $end
$var wire 1 #* c2 [16] $end
$var wire 1 $* c2 [15] $end
$var wire 1 %* c2 [14] $end
$var wire 1 &* c2 [13] $end
$var wire 1 '* c2 [12] $end
$var wire 1 (* c2 [11] $end
$var wire 1 )* c2 [10] $end
$var wire 1 ** c2 [9] $end
$var wire 1 +* c2 [8] $end
$var wire 1 ,* c2 [7] $end
$var wire 1 -* c2 [6] $end
$var wire 1 .* c2 [5] $end
$var wire 1 /* c2 [4] $end
$var wire 1 0* c2 [3] $end
$var wire 1 1* c2 [2] $end
$var wire 1 2* c2 [1] $end
$var wire 1 3* c2 [0] $end
$var wire 1 |* s [35] $end
$var wire 1 }* s [34] $end
$var wire 1 ~* s [33] $end
$var wire 1 !+ s [32] $end
$var wire 1 "+ s [31] $end
$var wire 1 #+ s [30] $end
$var wire 1 $+ s [29] $end
$var wire 1 %+ s [28] $end
$var wire 1 &+ s [27] $end
$var wire 1 '+ s [26] $end
$var wire 1 (+ s [25] $end
$var wire 1 )+ s [24] $end
$var wire 1 *+ s [23] $end
$var wire 1 ++ s [22] $end
$var wire 1 ,+ s [21] $end
$var wire 1 -+ s [20] $end
$var wire 1 .+ s [19] $end
$var wire 1 /+ s [18] $end
$var wire 1 0+ s [17] $end
$var wire 1 1+ s [16] $end
$var wire 1 2+ s [15] $end
$var wire 1 3+ s [14] $end
$var wire 1 4+ s [13] $end
$var wire 1 5+ s [12] $end
$var wire 1 6+ s [11] $end
$var wire 1 7+ s [10] $end
$var wire 1 8+ s [9] $end
$var wire 1 9+ s [8] $end
$var wire 1 :+ s [7] $end
$var wire 1 ;+ s [6] $end
$var wire 1 <+ s [5] $end
$var wire 1 =+ s [4] $end
$var wire 1 >+ s [3] $end
$var wire 1 ?+ s [2] $end
$var wire 1 @+ s [1] $end
$var wire 1 A+ s [0] $end
$var wire 1 B+ ca [35] $end
$var wire 1 C+ ca [34] $end
$var wire 1 D+ ca [33] $end
$var wire 1 E+ ca [32] $end
$var wire 1 F+ ca [31] $end
$var wire 1 G+ ca [30] $end
$var wire 1 H+ ca [29] $end
$var wire 1 I+ ca [28] $end
$var wire 1 J+ ca [27] $end
$var wire 1 K+ ca [26] $end
$var wire 1 L+ ca [25] $end
$var wire 1 M+ ca [24] $end
$var wire 1 N+ ca [23] $end
$var wire 1 O+ ca [22] $end
$var wire 1 P+ ca [21] $end
$var wire 1 Q+ ca [20] $end
$var wire 1 R+ ca [19] $end
$var wire 1 S+ ca [18] $end
$var wire 1 T+ ca [17] $end
$var wire 1 U+ ca [16] $end
$var wire 1 V+ ca [15] $end
$var wire 1 W+ ca [14] $end
$var wire 1 X+ ca [13] $end
$var wire 1 Y+ ca [12] $end
$var wire 1 Z+ ca [11] $end
$var wire 1 [+ ca [10] $end
$var wire 1 \+ ca [9] $end
$var wire 1 ]+ ca [8] $end
$var wire 1 ^+ ca [7] $end
$var wire 1 _+ ca [6] $end
$var wire 1 `+ ca [5] $end
$var wire 1 a+ ca [4] $end
$var wire 1 b+ ca [3] $end
$var wire 1 c+ ca [2] $end
$var wire 1 d+ ca [1] $end
$var wire 1 e+ ca [0] $end
$upscope $end

$scope module l1_2 $end
$var parameter 32 |Q size $end
$var wire 1 f+ c0 [39] $end
$var wire 1 g+ c0 [38] $end
$var wire 1 h+ c0 [37] $end
$var wire 1 i+ c0 [36] $end
$var wire 1 j+ c0 [35] $end
$var wire 1 k+ c0 [34] $end
$var wire 1 l+ c0 [33] $end
$var wire 1 m+ c0 [32] $end
$var wire 1 n+ c0 [31] $end
$var wire 1 o+ c0 [30] $end
$var wire 1 p+ c0 [29] $end
$var wire 1 q+ c0 [28] $end
$var wire 1 r+ c0 [27] $end
$var wire 1 s+ c0 [26] $end
$var wire 1 t+ c0 [25] $end
$var wire 1 u+ c0 [24] $end
$var wire 1 v+ c0 [23] $end
$var wire 1 w+ c0 [22] $end
$var wire 1 x+ c0 [21] $end
$var wire 1 y+ c0 [20] $end
$var wire 1 z+ c0 [19] $end
$var wire 1 {+ c0 [18] $end
$var wire 1 |+ c0 [17] $end
$var wire 1 }+ c0 [16] $end
$var wire 1 ~+ c0 [15] $end
$var wire 1 !, c0 [14] $end
$var wire 1 ", c0 [13] $end
$var wire 1 #, c0 [12] $end
$var wire 1 $, c0 [11] $end
$var wire 1 %, c0 [10] $end
$var wire 1 &, c0 [9] $end
$var wire 1 ', c0 [8] $end
$var wire 1 (, c0 [7] $end
$var wire 1 ), c0 [6] $end
$var wire 1 *, c0 [5] $end
$var wire 1 +, c0 [4] $end
$var wire 1 ,, c0 [3] $end
$var wire 1 -, c0 [2] $end
$var wire 1 ., c0 [1] $end
$var wire 1 /, c0 [0] $end
$var wire 1 0, c1 [39] $end
$var wire 1 1, c1 [38] $end
$var wire 1 2, c1 [37] $end
$var wire 1 3, c1 [36] $end
$var wire 1 4, c1 [35] $end
$var wire 1 5, c1 [34] $end
$var wire 1 6, c1 [33] $end
$var wire 1 7, c1 [32] $end
$var wire 1 8, c1 [31] $end
$var wire 1 9, c1 [30] $end
$var wire 1 :, c1 [29] $end
$var wire 1 ;, c1 [28] $end
$var wire 1 <, c1 [27] $end
$var wire 1 =, c1 [26] $end
$var wire 1 >, c1 [25] $end
$var wire 1 ?, c1 [24] $end
$var wire 1 @, c1 [23] $end
$var wire 1 A, c1 [22] $end
$var wire 1 B, c1 [21] $end
$var wire 1 C, c1 [20] $end
$var wire 1 D, c1 [19] $end
$var wire 1 E, c1 [18] $end
$var wire 1 F, c1 [17] $end
$var wire 1 G, c1 [16] $end
$var wire 1 H, c1 [15] $end
$var wire 1 I, c1 [14] $end
$var wire 1 J, c1 [13] $end
$var wire 1 K, c1 [12] $end
$var wire 1 L, c1 [11] $end
$var wire 1 M, c1 [10] $end
$var wire 1 N, c1 [9] $end
$var wire 1 O, c1 [8] $end
$var wire 1 P, c1 [7] $end
$var wire 1 Q, c1 [6] $end
$var wire 1 R, c1 [5] $end
$var wire 1 S, c1 [4] $end
$var wire 1 T, c1 [3] $end
$var wire 1 U, c1 [2] $end
$var wire 1 V, c1 [1] $end
$var wire 1 W, c1 [0] $end
$var wire 1 X, c2 [39] $end
$var wire 1 Y, c2 [38] $end
$var wire 1 Z, c2 [37] $end
$var wire 1 [, c2 [36] $end
$var wire 1 \, c2 [35] $end
$var wire 1 ], c2 [34] $end
$var wire 1 ^, c2 [33] $end
$var wire 1 _, c2 [32] $end
$var wire 1 `, c2 [31] $end
$var wire 1 a, c2 [30] $end
$var wire 1 b, c2 [29] $end
$var wire 1 c, c2 [28] $end
$var wire 1 d, c2 [27] $end
$var wire 1 e, c2 [26] $end
$var wire 1 f, c2 [25] $end
$var wire 1 g, c2 [24] $end
$var wire 1 h, c2 [23] $end
$var wire 1 i, c2 [22] $end
$var wire 1 j, c2 [21] $end
$var wire 1 k, c2 [20] $end
$var wire 1 l, c2 [19] $end
$var wire 1 m, c2 [18] $end
$var wire 1 n, c2 [17] $end
$var wire 1 o, c2 [16] $end
$var wire 1 p, c2 [15] $end
$var wire 1 q, c2 [14] $end
$var wire 1 r, c2 [13] $end
$var wire 1 s, c2 [12] $end
$var wire 1 t, c2 [11] $end
$var wire 1 u, c2 [10] $end
$var wire 1 v, c2 [9] $end
$var wire 1 w, c2 [8] $end
$var wire 1 x, c2 [7] $end
$var wire 1 y, c2 [6] $end
$var wire 1 z, c2 [5] $end
$var wire 1 {, c2 [4] $end
$var wire 1 |, c2 [3] $end
$var wire 1 }, c2 [2] $end
$var wire 1 ~, c2 [1] $end
$var wire 1 !- c2 [0] $end
$var wire 1 r- s [39] $end
$var wire 1 s- s [38] $end
$var wire 1 t- s [37] $end
$var wire 1 u- s [36] $end
$var wire 1 v- s [35] $end
$var wire 1 w- s [34] $end
$var wire 1 x- s [33] $end
$var wire 1 y- s [32] $end
$var wire 1 z- s [31] $end
$var wire 1 {- s [30] $end
$var wire 1 |- s [29] $end
$var wire 1 }- s [28] $end
$var wire 1 ~- s [27] $end
$var wire 1 !. s [26] $end
$var wire 1 ". s [25] $end
$var wire 1 #. s [24] $end
$var wire 1 $. s [23] $end
$var wire 1 %. s [22] $end
$var wire 1 &. s [21] $end
$var wire 1 '. s [20] $end
$var wire 1 (. s [19] $end
$var wire 1 ). s [18] $end
$var wire 1 *. s [17] $end
$var wire 1 +. s [16] $end
$var wire 1 ,. s [15] $end
$var wire 1 -. s [14] $end
$var wire 1 .. s [13] $end
$var wire 1 /. s [12] $end
$var wire 1 0. s [11] $end
$var wire 1 1. s [10] $end
$var wire 1 2. s [9] $end
$var wire 1 3. s [8] $end
$var wire 1 4. s [7] $end
$var wire 1 5. s [6] $end
$var wire 1 6. s [5] $end
$var wire 1 7. s [4] $end
$var wire 1 8. s [3] $end
$var wire 1 9. s [2] $end
$var wire 1 :. s [1] $end
$var wire 1 ;. s [0] $end
$var wire 1 <. ca [39] $end
$var wire 1 =. ca [38] $end
$var wire 1 >. ca [37] $end
$var wire 1 ?. ca [36] $end
$var wire 1 @. ca [35] $end
$var wire 1 A. ca [34] $end
$var wire 1 B. ca [33] $end
$var wire 1 C. ca [32] $end
$var wire 1 D. ca [31] $end
$var wire 1 E. ca [30] $end
$var wire 1 F. ca [29] $end
$var wire 1 G. ca [28] $end
$var wire 1 H. ca [27] $end
$var wire 1 I. ca [26] $end
$var wire 1 J. ca [25] $end
$var wire 1 K. ca [24] $end
$var wire 1 L. ca [23] $end
$var wire 1 M. ca [22] $end
$var wire 1 N. ca [21] $end
$var wire 1 O. ca [20] $end
$var wire 1 P. ca [19] $end
$var wire 1 Q. ca [18] $end
$var wire 1 R. ca [17] $end
$var wire 1 S. ca [16] $end
$var wire 1 T. ca [15] $end
$var wire 1 U. ca [14] $end
$var wire 1 V. ca [13] $end
$var wire 1 W. ca [12] $end
$var wire 1 X. ca [11] $end
$var wire 1 Y. ca [10] $end
$var wire 1 Z. ca [9] $end
$var wire 1 [. ca [8] $end
$var wire 1 \. ca [7] $end
$var wire 1 ]. ca [6] $end
$var wire 1 ^. ca [5] $end
$var wire 1 _. ca [4] $end
$var wire 1 `. ca [3] $end
$var wire 1 a. ca [2] $end
$var wire 1 b. ca [1] $end
$var wire 1 c. ca [0] $end
$upscope $end

$scope module l1_3 $end
$var parameter 32 }Q size $end
$var wire 1 d. c0 [39] $end
$var wire 1 e. c0 [38] $end
$var wire 1 f. c0 [37] $end
$var wire 1 g. c0 [36] $end
$var wire 1 h. c0 [35] $end
$var wire 1 i. c0 [34] $end
$var wire 1 j. c0 [33] $end
$var wire 1 k. c0 [32] $end
$var wire 1 l. c0 [31] $end
$var wire 1 m. c0 [30] $end
$var wire 1 n. c0 [29] $end
$var wire 1 o. c0 [28] $end
$var wire 1 p. c0 [27] $end
$var wire 1 q. c0 [26] $end
$var wire 1 r. c0 [25] $end
$var wire 1 s. c0 [24] $end
$var wire 1 t. c0 [23] $end
$var wire 1 u. c0 [22] $end
$var wire 1 v. c0 [21] $end
$var wire 1 w. c0 [20] $end
$var wire 1 x. c0 [19] $end
$var wire 1 y. c0 [18] $end
$var wire 1 z. c0 [17] $end
$var wire 1 {. c0 [16] $end
$var wire 1 |. c0 [15] $end
$var wire 1 }. c0 [14] $end
$var wire 1 ~. c0 [13] $end
$var wire 1 !/ c0 [12] $end
$var wire 1 "/ c0 [11] $end
$var wire 1 #/ c0 [10] $end
$var wire 1 $/ c0 [9] $end
$var wire 1 %/ c0 [8] $end
$var wire 1 &/ c0 [7] $end
$var wire 1 '/ c0 [6] $end
$var wire 1 (/ c0 [5] $end
$var wire 1 )/ c0 [4] $end
$var wire 1 */ c0 [3] $end
$var wire 1 +/ c0 [2] $end
$var wire 1 ,/ c0 [1] $end
$var wire 1 -/ c0 [0] $end
$var wire 1 ./ c1 [39] $end
$var wire 1 // c1 [38] $end
$var wire 1 0/ c1 [37] $end
$var wire 1 1/ c1 [36] $end
$var wire 1 2/ c1 [35] $end
$var wire 1 3/ c1 [34] $end
$var wire 1 4/ c1 [33] $end
$var wire 1 5/ c1 [32] $end
$var wire 1 6/ c1 [31] $end
$var wire 1 7/ c1 [30] $end
$var wire 1 8/ c1 [29] $end
$var wire 1 9/ c1 [28] $end
$var wire 1 :/ c1 [27] $end
$var wire 1 ;/ c1 [26] $end
$var wire 1 </ c1 [25] $end
$var wire 1 =/ c1 [24] $end
$var wire 1 >/ c1 [23] $end
$var wire 1 ?/ c1 [22] $end
$var wire 1 @/ c1 [21] $end
$var wire 1 A/ c1 [20] $end
$var wire 1 B/ c1 [19] $end
$var wire 1 C/ c1 [18] $end
$var wire 1 D/ c1 [17] $end
$var wire 1 E/ c1 [16] $end
$var wire 1 F/ c1 [15] $end
$var wire 1 G/ c1 [14] $end
$var wire 1 H/ c1 [13] $end
$var wire 1 I/ c1 [12] $end
$var wire 1 J/ c1 [11] $end
$var wire 1 K/ c1 [10] $end
$var wire 1 L/ c1 [9] $end
$var wire 1 M/ c1 [8] $end
$var wire 1 N/ c1 [7] $end
$var wire 1 O/ c1 [6] $end
$var wire 1 P/ c1 [5] $end
$var wire 1 Q/ c1 [4] $end
$var wire 1 R/ c1 [3] $end
$var wire 1 S/ c1 [2] $end
$var wire 1 T/ c1 [1] $end
$var wire 1 U/ c1 [0] $end
$var wire 1 V/ c2 [39] $end
$var wire 1 W/ c2 [38] $end
$var wire 1 X/ c2 [37] $end
$var wire 1 Y/ c2 [36] $end
$var wire 1 Z/ c2 [35] $end
$var wire 1 [/ c2 [34] $end
$var wire 1 \/ c2 [33] $end
$var wire 1 ]/ c2 [32] $end
$var wire 1 ^/ c2 [31] $end
$var wire 1 _/ c2 [30] $end
$var wire 1 `/ c2 [29] $end
$var wire 1 a/ c2 [28] $end
$var wire 1 b/ c2 [27] $end
$var wire 1 c/ c2 [26] $end
$var wire 1 d/ c2 [25] $end
$var wire 1 e/ c2 [24] $end
$var wire 1 f/ c2 [23] $end
$var wire 1 g/ c2 [22] $end
$var wire 1 h/ c2 [21] $end
$var wire 1 i/ c2 [20] $end
$var wire 1 j/ c2 [19] $end
$var wire 1 k/ c2 [18] $end
$var wire 1 l/ c2 [17] $end
$var wire 1 m/ c2 [16] $end
$var wire 1 n/ c2 [15] $end
$var wire 1 o/ c2 [14] $end
$var wire 1 p/ c2 [13] $end
$var wire 1 q/ c2 [12] $end
$var wire 1 r/ c2 [11] $end
$var wire 1 s/ c2 [10] $end
$var wire 1 t/ c2 [9] $end
$var wire 1 u/ c2 [8] $end
$var wire 1 v/ c2 [7] $end
$var wire 1 w/ c2 [6] $end
$var wire 1 x/ c2 [5] $end
$var wire 1 y/ c2 [4] $end
$var wire 1 z/ c2 [3] $end
$var wire 1 {/ c2 [2] $end
$var wire 1 |/ c2 [1] $end
$var wire 1 }/ c2 [0] $end
$var wire 1 p0 s [39] $end
$var wire 1 q0 s [38] $end
$var wire 1 r0 s [37] $end
$var wire 1 s0 s [36] $end
$var wire 1 t0 s [35] $end
$var wire 1 u0 s [34] $end
$var wire 1 v0 s [33] $end
$var wire 1 w0 s [32] $end
$var wire 1 x0 s [31] $end
$var wire 1 y0 s [30] $end
$var wire 1 z0 s [29] $end
$var wire 1 {0 s [28] $end
$var wire 1 |0 s [27] $end
$var wire 1 }0 s [26] $end
$var wire 1 ~0 s [25] $end
$var wire 1 !1 s [24] $end
$var wire 1 "1 s [23] $end
$var wire 1 #1 s [22] $end
$var wire 1 $1 s [21] $end
$var wire 1 %1 s [20] $end
$var wire 1 &1 s [19] $end
$var wire 1 '1 s [18] $end
$var wire 1 (1 s [17] $end
$var wire 1 )1 s [16] $end
$var wire 1 *1 s [15] $end
$var wire 1 +1 s [14] $end
$var wire 1 ,1 s [13] $end
$var wire 1 -1 s [12] $end
$var wire 1 .1 s [11] $end
$var wire 1 /1 s [10] $end
$var wire 1 01 s [9] $end
$var wire 1 11 s [8] $end
$var wire 1 21 s [7] $end
$var wire 1 31 s [6] $end
$var wire 1 41 s [5] $end
$var wire 1 51 s [4] $end
$var wire 1 61 s [3] $end
$var wire 1 71 s [2] $end
$var wire 1 81 s [1] $end
$var wire 1 91 s [0] $end
$var wire 1 :1 ca [39] $end
$var wire 1 ;1 ca [38] $end
$var wire 1 <1 ca [37] $end
$var wire 1 =1 ca [36] $end
$var wire 1 >1 ca [35] $end
$var wire 1 ?1 ca [34] $end
$var wire 1 @1 ca [33] $end
$var wire 1 A1 ca [32] $end
$var wire 1 B1 ca [31] $end
$var wire 1 C1 ca [30] $end
$var wire 1 D1 ca [29] $end
$var wire 1 E1 ca [28] $end
$var wire 1 F1 ca [27] $end
$var wire 1 G1 ca [26] $end
$var wire 1 H1 ca [25] $end
$var wire 1 I1 ca [24] $end
$var wire 1 J1 ca [23] $end
$var wire 1 K1 ca [22] $end
$var wire 1 L1 ca [21] $end
$var wire 1 M1 ca [20] $end
$var wire 1 N1 ca [19] $end
$var wire 1 O1 ca [18] $end
$var wire 1 P1 ca [17] $end
$var wire 1 Q1 ca [16] $end
$var wire 1 R1 ca [15] $end
$var wire 1 S1 ca [14] $end
$var wire 1 T1 ca [13] $end
$var wire 1 U1 ca [12] $end
$var wire 1 V1 ca [11] $end
$var wire 1 W1 ca [10] $end
$var wire 1 X1 ca [9] $end
$var wire 1 Y1 ca [8] $end
$var wire 1 Z1 ca [7] $end
$var wire 1 [1 ca [6] $end
$var wire 1 \1 ca [5] $end
$var wire 1 ]1 ca [4] $end
$var wire 1 ^1 ca [3] $end
$var wire 1 _1 ca [2] $end
$var wire 1 `1 ca [1] $end
$var wire 1 a1 ca [0] $end
$upscope $end

$scope module l1_4 $end
$var parameter 32 ~Q size $end
$var wire 1 b1 c0 [39] $end
$var wire 1 c1 c0 [38] $end
$var wire 1 d1 c0 [37] $end
$var wire 1 e1 c0 [36] $end
$var wire 1 f1 c0 [35] $end
$var wire 1 g1 c0 [34] $end
$var wire 1 h1 c0 [33] $end
$var wire 1 i1 c0 [32] $end
$var wire 1 j1 c0 [31] $end
$var wire 1 k1 c0 [30] $end
$var wire 1 l1 c0 [29] $end
$var wire 1 m1 c0 [28] $end
$var wire 1 n1 c0 [27] $end
$var wire 1 o1 c0 [26] $end
$var wire 1 p1 c0 [25] $end
$var wire 1 q1 c0 [24] $end
$var wire 1 r1 c0 [23] $end
$var wire 1 s1 c0 [22] $end
$var wire 1 t1 c0 [21] $end
$var wire 1 u1 c0 [20] $end
$var wire 1 v1 c0 [19] $end
$var wire 1 w1 c0 [18] $end
$var wire 1 x1 c0 [17] $end
$var wire 1 y1 c0 [16] $end
$var wire 1 z1 c0 [15] $end
$var wire 1 {1 c0 [14] $end
$var wire 1 |1 c0 [13] $end
$var wire 1 }1 c0 [12] $end
$var wire 1 ~1 c0 [11] $end
$var wire 1 !2 c0 [10] $end
$var wire 1 "2 c0 [9] $end
$var wire 1 #2 c0 [8] $end
$var wire 1 $2 c0 [7] $end
$var wire 1 %2 c0 [6] $end
$var wire 1 &2 c0 [5] $end
$var wire 1 '2 c0 [4] $end
$var wire 1 (2 c0 [3] $end
$var wire 1 )2 c0 [2] $end
$var wire 1 *2 c0 [1] $end
$var wire 1 +2 c0 [0] $end
$var wire 1 ,2 c1 [39] $end
$var wire 1 -2 c1 [38] $end
$var wire 1 .2 c1 [37] $end
$var wire 1 /2 c1 [36] $end
$var wire 1 02 c1 [35] $end
$var wire 1 12 c1 [34] $end
$var wire 1 22 c1 [33] $end
$var wire 1 32 c1 [32] $end
$var wire 1 42 c1 [31] $end
$var wire 1 52 c1 [30] $end
$var wire 1 62 c1 [29] $end
$var wire 1 72 c1 [28] $end
$var wire 1 82 c1 [27] $end
$var wire 1 92 c1 [26] $end
$var wire 1 :2 c1 [25] $end
$var wire 1 ;2 c1 [24] $end
$var wire 1 <2 c1 [23] $end
$var wire 1 =2 c1 [22] $end
$var wire 1 >2 c1 [21] $end
$var wire 1 ?2 c1 [20] $end
$var wire 1 @2 c1 [19] $end
$var wire 1 A2 c1 [18] $end
$var wire 1 B2 c1 [17] $end
$var wire 1 C2 c1 [16] $end
$var wire 1 D2 c1 [15] $end
$var wire 1 E2 c1 [14] $end
$var wire 1 F2 c1 [13] $end
$var wire 1 G2 c1 [12] $end
$var wire 1 H2 c1 [11] $end
$var wire 1 I2 c1 [10] $end
$var wire 1 J2 c1 [9] $end
$var wire 1 K2 c1 [8] $end
$var wire 1 L2 c1 [7] $end
$var wire 1 M2 c1 [6] $end
$var wire 1 N2 c1 [5] $end
$var wire 1 O2 c1 [4] $end
$var wire 1 P2 c1 [3] $end
$var wire 1 Q2 c1 [2] $end
$var wire 1 R2 c1 [1] $end
$var wire 1 S2 c1 [0] $end
$var wire 1 T2 c2 [39] $end
$var wire 1 U2 c2 [38] $end
$var wire 1 V2 c2 [37] $end
$var wire 1 W2 c2 [36] $end
$var wire 1 X2 c2 [35] $end
$var wire 1 Y2 c2 [34] $end
$var wire 1 Z2 c2 [33] $end
$var wire 1 [2 c2 [32] $end
$var wire 1 \2 c2 [31] $end
$var wire 1 ]2 c2 [30] $end
$var wire 1 ^2 c2 [29] $end
$var wire 1 _2 c2 [28] $end
$var wire 1 `2 c2 [27] $end
$var wire 1 a2 c2 [26] $end
$var wire 1 b2 c2 [25] $end
$var wire 1 c2 c2 [24] $end
$var wire 1 d2 c2 [23] $end
$var wire 1 e2 c2 [22] $end
$var wire 1 f2 c2 [21] $end
$var wire 1 g2 c2 [20] $end
$var wire 1 h2 c2 [19] $end
$var wire 1 i2 c2 [18] $end
$var wire 1 j2 c2 [17] $end
$var wire 1 k2 c2 [16] $end
$var wire 1 l2 c2 [15] $end
$var wire 1 m2 c2 [14] $end
$var wire 1 n2 c2 [13] $end
$var wire 1 o2 c2 [12] $end
$var wire 1 p2 c2 [11] $end
$var wire 1 q2 c2 [10] $end
$var wire 1 r2 c2 [9] $end
$var wire 1 s2 c2 [8] $end
$var wire 1 t2 c2 [7] $end
$var wire 1 u2 c2 [6] $end
$var wire 1 v2 c2 [5] $end
$var wire 1 w2 c2 [4] $end
$var wire 1 x2 c2 [3] $end
$var wire 1 y2 c2 [2] $end
$var wire 1 z2 c2 [1] $end
$var wire 1 {2 c2 [0] $end
$var wire 1 n3 s [39] $end
$var wire 1 o3 s [38] $end
$var wire 1 p3 s [37] $end
$var wire 1 q3 s [36] $end
$var wire 1 r3 s [35] $end
$var wire 1 s3 s [34] $end
$var wire 1 t3 s [33] $end
$var wire 1 u3 s [32] $end
$var wire 1 v3 s [31] $end
$var wire 1 w3 s [30] $end
$var wire 1 x3 s [29] $end
$var wire 1 y3 s [28] $end
$var wire 1 z3 s [27] $end
$var wire 1 {3 s [26] $end
$var wire 1 |3 s [25] $end
$var wire 1 }3 s [24] $end
$var wire 1 ~3 s [23] $end
$var wire 1 !4 s [22] $end
$var wire 1 "4 s [21] $end
$var wire 1 #4 s [20] $end
$var wire 1 $4 s [19] $end
$var wire 1 %4 s [18] $end
$var wire 1 &4 s [17] $end
$var wire 1 '4 s [16] $end
$var wire 1 (4 s [15] $end
$var wire 1 )4 s [14] $end
$var wire 1 *4 s [13] $end
$var wire 1 +4 s [12] $end
$var wire 1 ,4 s [11] $end
$var wire 1 -4 s [10] $end
$var wire 1 .4 s [9] $end
$var wire 1 /4 s [8] $end
$var wire 1 04 s [7] $end
$var wire 1 14 s [6] $end
$var wire 1 24 s [5] $end
$var wire 1 34 s [4] $end
$var wire 1 44 s [3] $end
$var wire 1 54 s [2] $end
$var wire 1 64 s [1] $end
$var wire 1 74 s [0] $end
$var wire 1 84 ca [39] $end
$var wire 1 94 ca [38] $end
$var wire 1 :4 ca [37] $end
$var wire 1 ;4 ca [36] $end
$var wire 1 <4 ca [35] $end
$var wire 1 =4 ca [34] $end
$var wire 1 >4 ca [33] $end
$var wire 1 ?4 ca [32] $end
$var wire 1 @4 ca [31] $end
$var wire 1 A4 ca [30] $end
$var wire 1 B4 ca [29] $end
$var wire 1 C4 ca [28] $end
$var wire 1 D4 ca [27] $end
$var wire 1 E4 ca [26] $end
$var wire 1 F4 ca [25] $end
$var wire 1 G4 ca [24] $end
$var wire 1 H4 ca [23] $end
$var wire 1 I4 ca [22] $end
$var wire 1 J4 ca [21] $end
$var wire 1 K4 ca [20] $end
$var wire 1 L4 ca [19] $end
$var wire 1 M4 ca [18] $end
$var wire 1 N4 ca [17] $end
$var wire 1 O4 ca [16] $end
$var wire 1 P4 ca [15] $end
$var wire 1 Q4 ca [14] $end
$var wire 1 R4 ca [13] $end
$var wire 1 S4 ca [12] $end
$var wire 1 T4 ca [11] $end
$var wire 1 U4 ca [10] $end
$var wire 1 V4 ca [9] $end
$var wire 1 W4 ca [8] $end
$var wire 1 X4 ca [7] $end
$var wire 1 Y4 ca [6] $end
$var wire 1 Z4 ca [5] $end
$var wire 1 [4 ca [4] $end
$var wire 1 \4 ca [3] $end
$var wire 1 ]4 ca [2] $end
$var wire 1 ^4 ca [1] $end
$var wire 1 _4 ca [0] $end
$upscope $end

$scope module l1_5 $end
$var parameter 32 !R size $end
$var wire 1 `4 c0 [39] $end
$var wire 1 a4 c0 [38] $end
$var wire 1 b4 c0 [37] $end
$var wire 1 c4 c0 [36] $end
$var wire 1 d4 c0 [35] $end
$var wire 1 e4 c0 [34] $end
$var wire 1 f4 c0 [33] $end
$var wire 1 g4 c0 [32] $end
$var wire 1 h4 c0 [31] $end
$var wire 1 i4 c0 [30] $end
$var wire 1 j4 c0 [29] $end
$var wire 1 k4 c0 [28] $end
$var wire 1 l4 c0 [27] $end
$var wire 1 m4 c0 [26] $end
$var wire 1 n4 c0 [25] $end
$var wire 1 o4 c0 [24] $end
$var wire 1 p4 c0 [23] $end
$var wire 1 q4 c0 [22] $end
$var wire 1 r4 c0 [21] $end
$var wire 1 s4 c0 [20] $end
$var wire 1 t4 c0 [19] $end
$var wire 1 u4 c0 [18] $end
$var wire 1 v4 c0 [17] $end
$var wire 1 w4 c0 [16] $end
$var wire 1 x4 c0 [15] $end
$var wire 1 y4 c0 [14] $end
$var wire 1 z4 c0 [13] $end
$var wire 1 {4 c0 [12] $end
$var wire 1 |4 c0 [11] $end
$var wire 1 }4 c0 [10] $end
$var wire 1 ~4 c0 [9] $end
$var wire 1 !5 c0 [8] $end
$var wire 1 "5 c0 [7] $end
$var wire 1 #5 c0 [6] $end
$var wire 1 $5 c0 [5] $end
$var wire 1 %5 c0 [4] $end
$var wire 1 &5 c0 [3] $end
$var wire 1 '5 c0 [2] $end
$var wire 1 (5 c0 [1] $end
$var wire 1 )5 c0 [0] $end
$var wire 1 *5 c1 [39] $end
$var wire 1 +5 c1 [38] $end
$var wire 1 ,5 c1 [37] $end
$var wire 1 -5 c1 [36] $end
$var wire 1 .5 c1 [35] $end
$var wire 1 /5 c1 [34] $end
$var wire 1 05 c1 [33] $end
$var wire 1 15 c1 [32] $end
$var wire 1 25 c1 [31] $end
$var wire 1 35 c1 [30] $end
$var wire 1 45 c1 [29] $end
$var wire 1 55 c1 [28] $end
$var wire 1 65 c1 [27] $end
$var wire 1 75 c1 [26] $end
$var wire 1 85 c1 [25] $end
$var wire 1 95 c1 [24] $end
$var wire 1 :5 c1 [23] $end
$var wire 1 ;5 c1 [22] $end
$var wire 1 <5 c1 [21] $end
$var wire 1 =5 c1 [20] $end
$var wire 1 >5 c1 [19] $end
$var wire 1 ?5 c1 [18] $end
$var wire 1 @5 c1 [17] $end
$var wire 1 A5 c1 [16] $end
$var wire 1 B5 c1 [15] $end
$var wire 1 C5 c1 [14] $end
$var wire 1 D5 c1 [13] $end
$var wire 1 E5 c1 [12] $end
$var wire 1 F5 c1 [11] $end
$var wire 1 G5 c1 [10] $end
$var wire 1 H5 c1 [9] $end
$var wire 1 I5 c1 [8] $end
$var wire 1 J5 c1 [7] $end
$var wire 1 K5 c1 [6] $end
$var wire 1 L5 c1 [5] $end
$var wire 1 M5 c1 [4] $end
$var wire 1 N5 c1 [3] $end
$var wire 1 O5 c1 [2] $end
$var wire 1 P5 c1 [1] $end
$var wire 1 Q5 c1 [0] $end
$var wire 1 R5 c2 [39] $end
$var wire 1 S5 c2 [38] $end
$var wire 1 T5 c2 [37] $end
$var wire 1 U5 c2 [36] $end
$var wire 1 V5 c2 [35] $end
$var wire 1 W5 c2 [34] $end
$var wire 1 X5 c2 [33] $end
$var wire 1 Y5 c2 [32] $end
$var wire 1 Z5 c2 [31] $end
$var wire 1 [5 c2 [30] $end
$var wire 1 \5 c2 [29] $end
$var wire 1 ]5 c2 [28] $end
$var wire 1 ^5 c2 [27] $end
$var wire 1 _5 c2 [26] $end
$var wire 1 `5 c2 [25] $end
$var wire 1 a5 c2 [24] $end
$var wire 1 b5 c2 [23] $end
$var wire 1 c5 c2 [22] $end
$var wire 1 d5 c2 [21] $end
$var wire 1 e5 c2 [20] $end
$var wire 1 f5 c2 [19] $end
$var wire 1 g5 c2 [18] $end
$var wire 1 h5 c2 [17] $end
$var wire 1 i5 c2 [16] $end
$var wire 1 j5 c2 [15] $end
$var wire 1 k5 c2 [14] $end
$var wire 1 l5 c2 [13] $end
$var wire 1 m5 c2 [12] $end
$var wire 1 n5 c2 [11] $end
$var wire 1 o5 c2 [10] $end
$var wire 1 p5 c2 [9] $end
$var wire 1 q5 c2 [8] $end
$var wire 1 r5 c2 [7] $end
$var wire 1 s5 c2 [6] $end
$var wire 1 t5 c2 [5] $end
$var wire 1 u5 c2 [4] $end
$var wire 1 v5 c2 [3] $end
$var wire 1 w5 c2 [2] $end
$var wire 1 x5 c2 [1] $end
$var wire 1 y5 c2 [0] $end
$var wire 1 l6 s [39] $end
$var wire 1 m6 s [38] $end
$var wire 1 n6 s [37] $end
$var wire 1 o6 s [36] $end
$var wire 1 p6 s [35] $end
$var wire 1 q6 s [34] $end
$var wire 1 r6 s [33] $end
$var wire 1 s6 s [32] $end
$var wire 1 t6 s [31] $end
$var wire 1 u6 s [30] $end
$var wire 1 v6 s [29] $end
$var wire 1 w6 s [28] $end
$var wire 1 x6 s [27] $end
$var wire 1 y6 s [26] $end
$var wire 1 z6 s [25] $end
$var wire 1 {6 s [24] $end
$var wire 1 |6 s [23] $end
$var wire 1 }6 s [22] $end
$var wire 1 ~6 s [21] $end
$var wire 1 !7 s [20] $end
$var wire 1 "7 s [19] $end
$var wire 1 #7 s [18] $end
$var wire 1 $7 s [17] $end
$var wire 1 %7 s [16] $end
$var wire 1 &7 s [15] $end
$var wire 1 '7 s [14] $end
$var wire 1 (7 s [13] $end
$var wire 1 )7 s [12] $end
$var wire 1 *7 s [11] $end
$var wire 1 +7 s [10] $end
$var wire 1 ,7 s [9] $end
$var wire 1 -7 s [8] $end
$var wire 1 .7 s [7] $end
$var wire 1 /7 s [6] $end
$var wire 1 07 s [5] $end
$var wire 1 17 s [4] $end
$var wire 1 27 s [3] $end
$var wire 1 37 s [2] $end
$var wire 1 47 s [1] $end
$var wire 1 57 s [0] $end
$var wire 1 67 ca [39] $end
$var wire 1 77 ca [38] $end
$var wire 1 87 ca [37] $end
$var wire 1 97 ca [36] $end
$var wire 1 :7 ca [35] $end
$var wire 1 ;7 ca [34] $end
$var wire 1 <7 ca [33] $end
$var wire 1 =7 ca [32] $end
$var wire 1 >7 ca [31] $end
$var wire 1 ?7 ca [30] $end
$var wire 1 @7 ca [29] $end
$var wire 1 A7 ca [28] $end
$var wire 1 B7 ca [27] $end
$var wire 1 C7 ca [26] $end
$var wire 1 D7 ca [25] $end
$var wire 1 E7 ca [24] $end
$var wire 1 F7 ca [23] $end
$var wire 1 G7 ca [22] $end
$var wire 1 H7 ca [21] $end
$var wire 1 I7 ca [20] $end
$var wire 1 J7 ca [19] $end
$var wire 1 K7 ca [18] $end
$var wire 1 L7 ca [17] $end
$var wire 1 M7 ca [16] $end
$var wire 1 N7 ca [15] $end
$var wire 1 O7 ca [14] $end
$var wire 1 P7 ca [13] $end
$var wire 1 Q7 ca [12] $end
$var wire 1 R7 ca [11] $end
$var wire 1 S7 ca [10] $end
$var wire 1 T7 ca [9] $end
$var wire 1 U7 ca [8] $end
$var wire 1 V7 ca [7] $end
$var wire 1 W7 ca [6] $end
$var wire 1 X7 ca [5] $end
$var wire 1 Y7 ca [4] $end
$var wire 1 Z7 ca [3] $end
$var wire 1 [7 ca [2] $end
$var wire 1 \7 ca [1] $end
$var wire 1 ]7 ca [0] $end
$upscope $end

$scope module l1_6 $end
$var parameter 32 "R size $end
$var wire 1 ^7 c0 [37] $end
$var wire 1 _7 c0 [36] $end
$var wire 1 `7 c0 [35] $end
$var wire 1 a7 c0 [34] $end
$var wire 1 b7 c0 [33] $end
$var wire 1 c7 c0 [32] $end
$var wire 1 d7 c0 [31] $end
$var wire 1 e7 c0 [30] $end
$var wire 1 f7 c0 [29] $end
$var wire 1 g7 c0 [28] $end
$var wire 1 h7 c0 [27] $end
$var wire 1 i7 c0 [26] $end
$var wire 1 j7 c0 [25] $end
$var wire 1 k7 c0 [24] $end
$var wire 1 l7 c0 [23] $end
$var wire 1 m7 c0 [22] $end
$var wire 1 n7 c0 [21] $end
$var wire 1 o7 c0 [20] $end
$var wire 1 p7 c0 [19] $end
$var wire 1 q7 c0 [18] $end
$var wire 1 r7 c0 [17] $end
$var wire 1 s7 c0 [16] $end
$var wire 1 t7 c0 [15] $end
$var wire 1 u7 c0 [14] $end
$var wire 1 v7 c0 [13] $end
$var wire 1 w7 c0 [12] $end
$var wire 1 x7 c0 [11] $end
$var wire 1 y7 c0 [10] $end
$var wire 1 z7 c0 [9] $end
$var wire 1 {7 c0 [8] $end
$var wire 1 |7 c0 [7] $end
$var wire 1 }7 c0 [6] $end
$var wire 1 ~7 c0 [5] $end
$var wire 1 !8 c0 [4] $end
$var wire 1 "8 c0 [3] $end
$var wire 1 #8 c0 [2] $end
$var wire 1 $8 c0 [1] $end
$var wire 1 %8 c0 [0] $end
$var wire 1 &8 c1 [37] $end
$var wire 1 '8 c1 [36] $end
$var wire 1 (8 c1 [35] $end
$var wire 1 )8 c1 [34] $end
$var wire 1 *8 c1 [33] $end
$var wire 1 +8 c1 [32] $end
$var wire 1 ,8 c1 [31] $end
$var wire 1 -8 c1 [30] $end
$var wire 1 .8 c1 [29] $end
$var wire 1 /8 c1 [28] $end
$var wire 1 08 c1 [27] $end
$var wire 1 18 c1 [26] $end
$var wire 1 28 c1 [25] $end
$var wire 1 38 c1 [24] $end
$var wire 1 48 c1 [23] $end
$var wire 1 58 c1 [22] $end
$var wire 1 68 c1 [21] $end
$var wire 1 78 c1 [20] $end
$var wire 1 88 c1 [19] $end
$var wire 1 98 c1 [18] $end
$var wire 1 :8 c1 [17] $end
$var wire 1 ;8 c1 [16] $end
$var wire 1 <8 c1 [15] $end
$var wire 1 =8 c1 [14] $end
$var wire 1 >8 c1 [13] $end
$var wire 1 ?8 c1 [12] $end
$var wire 1 @8 c1 [11] $end
$var wire 1 A8 c1 [10] $end
$var wire 1 B8 c1 [9] $end
$var wire 1 C8 c1 [8] $end
$var wire 1 D8 c1 [7] $end
$var wire 1 E8 c1 [6] $end
$var wire 1 F8 c1 [5] $end
$var wire 1 G8 c1 [4] $end
$var wire 1 H8 c1 [3] $end
$var wire 1 I8 c1 [2] $end
$var wire 1 J8 c1 [1] $end
$var wire 1 K8 c1 [0] $end
$var wire 1 L8 c2 [37] $end
$var wire 1 M8 c2 [36] $end
$var wire 1 N8 c2 [35] $end
$var wire 1 O8 c2 [34] $end
$var wire 1 P8 c2 [33] $end
$var wire 1 Q8 c2 [32] $end
$var wire 1 R8 c2 [31] $end
$var wire 1 S8 c2 [30] $end
$var wire 1 T8 c2 [29] $end
$var wire 1 U8 c2 [28] $end
$var wire 1 V8 c2 [27] $end
$var wire 1 W8 c2 [26] $end
$var wire 1 X8 c2 [25] $end
$var wire 1 Y8 c2 [24] $end
$var wire 1 Z8 c2 [23] $end
$var wire 1 [8 c2 [22] $end
$var wire 1 \8 c2 [21] $end
$var wire 1 ]8 c2 [20] $end
$var wire 1 ^8 c2 [19] $end
$var wire 1 _8 c2 [18] $end
$var wire 1 `8 c2 [17] $end
$var wire 1 a8 c2 [16] $end
$var wire 1 b8 c2 [15] $end
$var wire 1 c8 c2 [14] $end
$var wire 1 d8 c2 [13] $end
$var wire 1 e8 c2 [12] $end
$var wire 1 f8 c2 [11] $end
$var wire 1 g8 c2 [10] $end
$var wire 1 h8 c2 [9] $end
$var wire 1 i8 c2 [8] $end
$var wire 1 j8 c2 [7] $end
$var wire 1 k8 c2 [6] $end
$var wire 1 l8 c2 [5] $end
$var wire 1 m8 c2 [4] $end
$var wire 1 n8 c2 [3] $end
$var wire 1 o8 c2 [2] $end
$var wire 1 p8 c2 [1] $end
$var wire 1 q8 c2 [0] $end
$var wire 1 `9 s [37] $end
$var wire 1 a9 s [36] $end
$var wire 1 b9 s [35] $end
$var wire 1 c9 s [34] $end
$var wire 1 d9 s [33] $end
$var wire 1 e9 s [32] $end
$var wire 1 f9 s [31] $end
$var wire 1 g9 s [30] $end
$var wire 1 h9 s [29] $end
$var wire 1 i9 s [28] $end
$var wire 1 j9 s [27] $end
$var wire 1 k9 s [26] $end
$var wire 1 l9 s [25] $end
$var wire 1 m9 s [24] $end
$var wire 1 n9 s [23] $end
$var wire 1 o9 s [22] $end
$var wire 1 p9 s [21] $end
$var wire 1 q9 s [20] $end
$var wire 1 r9 s [19] $end
$var wire 1 s9 s [18] $end
$var wire 1 t9 s [17] $end
$var wire 1 u9 s [16] $end
$var wire 1 v9 s [15] $end
$var wire 1 w9 s [14] $end
$var wire 1 x9 s [13] $end
$var wire 1 y9 s [12] $end
$var wire 1 z9 s [11] $end
$var wire 1 {9 s [10] $end
$var wire 1 |9 s [9] $end
$var wire 1 }9 s [8] $end
$var wire 1 ~9 s [7] $end
$var wire 1 !: s [6] $end
$var wire 1 ": s [5] $end
$var wire 1 #: s [4] $end
$var wire 1 $: s [3] $end
$var wire 1 %: s [2] $end
$var wire 1 &: s [1] $end
$var wire 1 ': s [0] $end
$var wire 1 (: ca [37] $end
$var wire 1 ): ca [36] $end
$var wire 1 *: ca [35] $end
$var wire 1 +: ca [34] $end
$var wire 1 ,: ca [33] $end
$var wire 1 -: ca [32] $end
$var wire 1 .: ca [31] $end
$var wire 1 /: ca [30] $end
$var wire 1 0: ca [29] $end
$var wire 1 1: ca [28] $end
$var wire 1 2: ca [27] $end
$var wire 1 3: ca [26] $end
$var wire 1 4: ca [25] $end
$var wire 1 5: ca [24] $end
$var wire 1 6: ca [23] $end
$var wire 1 7: ca [22] $end
$var wire 1 8: ca [21] $end
$var wire 1 9: ca [20] $end
$var wire 1 :: ca [19] $end
$var wire 1 ;: ca [18] $end
$var wire 1 <: ca [17] $end
$var wire 1 =: ca [16] $end
$var wire 1 >: ca [15] $end
$var wire 1 ?: ca [14] $end
$var wire 1 @: ca [13] $end
$var wire 1 A: ca [12] $end
$var wire 1 B: ca [11] $end
$var wire 1 C: ca [10] $end
$var wire 1 D: ca [9] $end
$var wire 1 E: ca [8] $end
$var wire 1 F: ca [7] $end
$var wire 1 G: ca [6] $end
$var wire 1 H: ca [5] $end
$var wire 1 I: ca [4] $end
$var wire 1 J: ca [3] $end
$var wire 1 K: ca [2] $end
$var wire 1 L: ca [1] $end
$var wire 1 M: ca [0] $end
$upscope $end

$scope module l2_1 $end
$var parameter 32 #R size $end
$var wire 1 $R p1 [42] $end
$var wire 1 %R p1 [41] $end
$var wire 1 &R p1 [40] $end
$var wire 1 'R p1 [39] $end
$var wire 1 (R p1 [38] $end
$var wire 1 )R p1 [37] $end
$var wire 1 *R p1 [36] $end
$var wire 1 +R p1 [35] $end
$var wire 1 ,R p1 [34] $end
$var wire 1 -R p1 [33] $end
$var wire 1 .R p1 [32] $end
$var wire 1 /R p1 [31] $end
$var wire 1 0R p1 [30] $end
$var wire 1 1R p1 [29] $end
$var wire 1 2R p1 [28] $end
$var wire 1 3R p1 [27] $end
$var wire 1 4R p1 [26] $end
$var wire 1 5R p1 [25] $end
$var wire 1 6R p1 [24] $end
$var wire 1 7R p1 [23] $end
$var wire 1 8R p1 [22] $end
$var wire 1 9R p1 [21] $end
$var wire 1 :R p1 [20] $end
$var wire 1 ;R p1 [19] $end
$var wire 1 <R p1 [18] $end
$var wire 1 =R p1 [17] $end
$var wire 1 >R p1 [16] $end
$var wire 1 ?R p1 [15] $end
$var wire 1 @R p1 [14] $end
$var wire 1 AR p1 [13] $end
$var wire 1 BR p1 [12] $end
$var wire 1 CR p1 [11] $end
$var wire 1 DR p1 [10] $end
$var wire 1 ER p1 [9] $end
$var wire 1 FR p1 [8] $end
$var wire 1 GR p1 [7] $end
$var wire 1 HR p1 [6] $end
$var wire 1 IR p1 [5] $end
$var wire 1 JR p1 [4] $end
$var wire 1 KR p1 [3] $end
$var wire 1 LR p1 [2] $end
$var wire 1 MR p1 [1] $end
$var wire 1 NR p1 [0] $end
$var wire 1 OR p2 [42] $end
$var wire 1 PR p2 [41] $end
$var wire 1 QR p2 [40] $end
$var wire 1 RR p2 [39] $end
$var wire 1 SR p2 [38] $end
$var wire 1 TR p2 [37] $end
$var wire 1 UR p2 [36] $end
$var wire 1 VR p2 [35] $end
$var wire 1 WR p2 [34] $end
$var wire 1 XR p2 [33] $end
$var wire 1 YR p2 [32] $end
$var wire 1 ZR p2 [31] $end
$var wire 1 [R p2 [30] $end
$var wire 1 \R p2 [29] $end
$var wire 1 ]R p2 [28] $end
$var wire 1 ^R p2 [27] $end
$var wire 1 _R p2 [26] $end
$var wire 1 `R p2 [25] $end
$var wire 1 aR p2 [24] $end
$var wire 1 bR p2 [23] $end
$var wire 1 cR p2 [22] $end
$var wire 1 dR p2 [21] $end
$var wire 1 eR p2 [20] $end
$var wire 1 fR p2 [19] $end
$var wire 1 gR p2 [18] $end
$var wire 1 hR p2 [17] $end
$var wire 1 iR p2 [16] $end
$var wire 1 jR p2 [15] $end
$var wire 1 kR p2 [14] $end
$var wire 1 lR p2 [13] $end
$var wire 1 mR p2 [12] $end
$var wire 1 nR p2 [11] $end
$var wire 1 oR p2 [10] $end
$var wire 1 pR p2 [9] $end
$var wire 1 qR p2 [8] $end
$var wire 1 rR p2 [7] $end
$var wire 1 sR p2 [6] $end
$var wire 1 tR p2 [5] $end
$var wire 1 uR p2 [4] $end
$var wire 1 vR p2 [3] $end
$var wire 1 wR p2 [2] $end
$var wire 1 xR p2 [1] $end
$var wire 1 yR p2 [0] $end
$var wire 1 zR p3 [42] $end
$var wire 1 {R p3 [41] $end
$var wire 1 |R p3 [40] $end
$var wire 1 }R p3 [39] $end
$var wire 1 ~R p3 [38] $end
$var wire 1 !S p3 [37] $end
$var wire 1 "S p3 [36] $end
$var wire 1 #S p3 [35] $end
$var wire 1 $S p3 [34] $end
$var wire 1 %S p3 [33] $end
$var wire 1 &S p3 [32] $end
$var wire 1 'S p3 [31] $end
$var wire 1 (S p3 [30] $end
$var wire 1 )S p3 [29] $end
$var wire 1 *S p3 [28] $end
$var wire 1 +S p3 [27] $end
$var wire 1 ,S p3 [26] $end
$var wire 1 -S p3 [25] $end
$var wire 1 .S p3 [24] $end
$var wire 1 /S p3 [23] $end
$var wire 1 0S p3 [22] $end
$var wire 1 1S p3 [21] $end
$var wire 1 2S p3 [20] $end
$var wire 1 3S p3 [19] $end
$var wire 1 4S p3 [18] $end
$var wire 1 5S p3 [17] $end
$var wire 1 6S p3 [16] $end
$var wire 1 7S p3 [15] $end
$var wire 1 8S p3 [14] $end
$var wire 1 9S p3 [13] $end
$var wire 1 :S p3 [12] $end
$var wire 1 ;S p3 [11] $end
$var wire 1 <S p3 [10] $end
$var wire 1 =S p3 [9] $end
$var wire 1 >S p3 [8] $end
$var wire 1 ?S p3 [7] $end
$var wire 1 @S p3 [6] $end
$var wire 1 AS p3 [5] $end
$var wire 1 BS p3 [4] $end
$var wire 1 CS p3 [3] $end
$var wire 1 DS p3 [2] $end
$var wire 1 ES p3 [1] $end
$var wire 1 FS p3 [0] $end
$var wire 1 Z: c1 [42] $end
$var wire 1 [: c1 [41] $end
$var wire 1 \: c1 [40] $end
$var wire 1 ]: c1 [39] $end
$var wire 1 ^: c1 [38] $end
$var wire 1 _: c1 [37] $end
$var wire 1 `: c1 [36] $end
$var wire 1 a: c1 [35] $end
$var wire 1 b: c1 [34] $end
$var wire 1 c: c1 [33] $end
$var wire 1 d: c1 [32] $end
$var wire 1 e: c1 [31] $end
$var wire 1 f: c1 [30] $end
$var wire 1 g: c1 [29] $end
$var wire 1 h: c1 [28] $end
$var wire 1 i: c1 [27] $end
$var wire 1 j: c1 [26] $end
$var wire 1 k: c1 [25] $end
$var wire 1 l: c1 [24] $end
$var wire 1 m: c1 [23] $end
$var wire 1 n: c1 [22] $end
$var wire 1 o: c1 [21] $end
$var wire 1 p: c1 [20] $end
$var wire 1 q: c1 [19] $end
$var wire 1 r: c1 [18] $end
$var wire 1 s: c1 [17] $end
$var wire 1 t: c1 [16] $end
$var wire 1 u: c1 [15] $end
$var wire 1 v: c1 [14] $end
$var wire 1 w: c1 [13] $end
$var wire 1 x: c1 [12] $end
$var wire 1 y: c1 [11] $end
$var wire 1 z: c1 [10] $end
$var wire 1 {: c1 [9] $end
$var wire 1 |: c1 [8] $end
$var wire 1 }: c1 [7] $end
$var wire 1 ~: c1 [6] $end
$var wire 1 !; c1 [5] $end
$var wire 1 "; c1 [4] $end
$var wire 1 #; c1 [3] $end
$var wire 1 $; c1 [2] $end
$var wire 1 %; c1 [1] $end
$var wire 1 &; c1 [0] $end
$var wire 1 '; c2 [42] $end
$var wire 1 (; c2 [41] $end
$var wire 1 ); c2 [40] $end
$var wire 1 *; c2 [39] $end
$var wire 1 +; c2 [38] $end
$var wire 1 ,; c2 [37] $end
$var wire 1 -; c2 [36] $end
$var wire 1 .; c2 [35] $end
$var wire 1 /; c2 [34] $end
$var wire 1 0; c2 [33] $end
$var wire 1 1; c2 [32] $end
$var wire 1 2; c2 [31] $end
$var wire 1 3; c2 [30] $end
$var wire 1 4; c2 [29] $end
$var wire 1 5; c2 [28] $end
$var wire 1 6; c2 [27] $end
$var wire 1 7; c2 [26] $end
$var wire 1 8; c2 [25] $end
$var wire 1 9; c2 [24] $end
$var wire 1 :; c2 [23] $end
$var wire 1 ;; c2 [22] $end
$var wire 1 <; c2 [21] $end
$var wire 1 =; c2 [20] $end
$var wire 1 >; c2 [19] $end
$var wire 1 ?; c2 [18] $end
$var wire 1 @; c2 [17] $end
$var wire 1 A; c2 [16] $end
$var wire 1 B; c2 [15] $end
$var wire 1 C; c2 [14] $end
$var wire 1 D; c2 [13] $end
$var wire 1 E; c2 [12] $end
$var wire 1 F; c2 [11] $end
$var wire 1 G; c2 [10] $end
$var wire 1 H; c2 [9] $end
$var wire 1 I; c2 [8] $end
$var wire 1 J; c2 [7] $end
$var wire 1 K; c2 [6] $end
$var wire 1 L; c2 [5] $end
$var wire 1 M; c2 [4] $end
$var wire 1 N; c2 [3] $end
$var wire 1 O; c2 [2] $end
$var wire 1 P; c2 [1] $end
$var wire 1 Q; c2 [0] $end
$var wire 1 R; c3 [42] $end
$var wire 1 S; c3 [41] $end
$var wire 1 T; c3 [40] $end
$var wire 1 U; c3 [39] $end
$var wire 1 V; c3 [38] $end
$var wire 1 W; c3 [37] $end
$var wire 1 X; c3 [36] $end
$var wire 1 Y; c3 [35] $end
$var wire 1 Z; c3 [34] $end
$var wire 1 [; c3 [33] $end
$var wire 1 \; c3 [32] $end
$var wire 1 ]; c3 [31] $end
$var wire 1 ^; c3 [30] $end
$var wire 1 _; c3 [29] $end
$var wire 1 `; c3 [28] $end
$var wire 1 a; c3 [27] $end
$var wire 1 b; c3 [26] $end
$var wire 1 c; c3 [25] $end
$var wire 1 d; c3 [24] $end
$var wire 1 e; c3 [23] $end
$var wire 1 f; c3 [22] $end
$var wire 1 g; c3 [21] $end
$var wire 1 h; c3 [20] $end
$var wire 1 i; c3 [19] $end
$var wire 1 j; c3 [18] $end
$var wire 1 k; c3 [17] $end
$var wire 1 l; c3 [16] $end
$var wire 1 m; c3 [15] $end
$var wire 1 n; c3 [14] $end
$var wire 1 o; c3 [13] $end
$var wire 1 p; c3 [12] $end
$var wire 1 q; c3 [11] $end
$var wire 1 r; c3 [10] $end
$var wire 1 s; c3 [9] $end
$var wire 1 t; c3 [8] $end
$var wire 1 u; c3 [7] $end
$var wire 1 v; c3 [6] $end
$var wire 1 w; c3 [5] $end
$var wire 1 x; c3 [4] $end
$var wire 1 y; c3 [3] $end
$var wire 1 z; c3 [2] $end
$var wire 1 {; c3 [1] $end
$var wire 1 |; c3 [0] $end
$var wire 1 }; c4 [42] $end
$var wire 1 ~; c4 [41] $end
$var wire 1 !< c4 [40] $end
$var wire 1 "< c4 [39] $end
$var wire 1 #< c4 [38] $end
$var wire 1 $< c4 [37] $end
$var wire 1 %< c4 [36] $end
$var wire 1 &< c4 [35] $end
$var wire 1 '< c4 [34] $end
$var wire 1 (< c4 [33] $end
$var wire 1 )< c4 [32] $end
$var wire 1 *< c4 [31] $end
$var wire 1 +< c4 [30] $end
$var wire 1 ,< c4 [29] $end
$var wire 1 -< c4 [28] $end
$var wire 1 .< c4 [27] $end
$var wire 1 /< c4 [26] $end
$var wire 1 0< c4 [25] $end
$var wire 1 1< c4 [24] $end
$var wire 1 2< c4 [23] $end
$var wire 1 3< c4 [22] $end
$var wire 1 4< c4 [21] $end
$var wire 1 5< c4 [20] $end
$var wire 1 6< c4 [19] $end
$var wire 1 7< c4 [18] $end
$var wire 1 8< c4 [17] $end
$var wire 1 9< c4 [16] $end
$var wire 1 :< c4 [15] $end
$var wire 1 ;< c4 [14] $end
$var wire 1 << c4 [13] $end
$var wire 1 =< c4 [12] $end
$var wire 1 >< c4 [11] $end
$var wire 1 ?< c4 [10] $end
$var wire 1 @< c4 [9] $end
$var wire 1 A< c4 [8] $end
$var wire 1 B< c4 [7] $end
$var wire 1 C< c4 [6] $end
$var wire 1 D< c4 [5] $end
$var wire 1 E< c4 [4] $end
$var wire 1 F< c4 [3] $end
$var wire 1 G< c4 [2] $end
$var wire 1 H< c4 [1] $end
$var wire 1 I< c4 [0] $end
$var wire 1 J< cin [42] $end
$var wire 1 K< cin [41] $end
$var wire 1 L< cin [40] $end
$var wire 1 M< cin [39] $end
$var wire 1 N< cin [38] $end
$var wire 1 O< cin [37] $end
$var wire 1 P< cin [36] $end
$var wire 1 Q< cin [35] $end
$var wire 1 R< cin [34] $end
$var wire 1 S< cin [33] $end
$var wire 1 T< cin [32] $end
$var wire 1 U< cin [31] $end
$var wire 1 V< cin [30] $end
$var wire 1 W< cin [29] $end
$var wire 1 X< cin [28] $end
$var wire 1 Y< cin [27] $end
$var wire 1 Z< cin [26] $end
$var wire 1 [< cin [25] $end
$var wire 1 \< cin [24] $end
$var wire 1 ]< cin [23] $end
$var wire 1 ^< cin [22] $end
$var wire 1 _< cin [21] $end
$var wire 1 `< cin [20] $end
$var wire 1 a< cin [19] $end
$var wire 1 b< cin [18] $end
$var wire 1 c< cin [17] $end
$var wire 1 d< cin [16] $end
$var wire 1 e< cin [15] $end
$var wire 1 f< cin [14] $end
$var wire 1 g< cin [13] $end
$var wire 1 h< cin [12] $end
$var wire 1 i< cin [11] $end
$var wire 1 j< cin [10] $end
$var wire 1 k< cin [9] $end
$var wire 1 l< cin [8] $end
$var wire 1 m< cin [7] $end
$var wire 1 n< cin [6] $end
$var wire 1 o< cin [5] $end
$var wire 1 p< cin [4] $end
$var wire 1 q< cin [3] $end
$var wire 1 r< cin [2] $end
$var wire 1 s< cin [1] $end
$var wire 1 t< cin [0] $end
$var wire 1 u< cout [42] $end
$var wire 1 v< cout [41] $end
$var wire 1 w< cout [40] $end
$var wire 1 x< cout [39] $end
$var wire 1 y< cout [38] $end
$var wire 1 z< cout [37] $end
$var wire 1 {< cout [36] $end
$var wire 1 |< cout [35] $end
$var wire 1 }< cout [34] $end
$var wire 1 ~< cout [33] $end
$var wire 1 != cout [32] $end
$var wire 1 "= cout [31] $end
$var wire 1 #= cout [30] $end
$var wire 1 $= cout [29] $end
$var wire 1 %= cout [28] $end
$var wire 1 &= cout [27] $end
$var wire 1 '= cout [26] $end
$var wire 1 (= cout [25] $end
$var wire 1 )= cout [24] $end
$var wire 1 *= cout [23] $end
$var wire 1 += cout [22] $end
$var wire 1 ,= cout [21] $end
$var wire 1 -= cout [20] $end
$var wire 1 .= cout [19] $end
$var wire 1 /= cout [18] $end
$var wire 1 0= cout [17] $end
$var wire 1 1= cout [16] $end
$var wire 1 2= cout [15] $end
$var wire 1 3= cout [14] $end
$var wire 1 4= cout [13] $end
$var wire 1 5= cout [12] $end
$var wire 1 6= cout [11] $end
$var wire 1 7= cout [10] $end
$var wire 1 8= cout [9] $end
$var wire 1 9= cout [8] $end
$var wire 1 := cout [7] $end
$var wire 1 ;= cout [6] $end
$var wire 1 <= cout [5] $end
$var wire 1 == cout [4] $end
$var wire 1 >= cout [3] $end
$var wire 1 ?= cout [2] $end
$var wire 1 @= cout [1] $end
$var wire 1 A= cout [0] $end
$var wire 1 B= s [42] $end
$var wire 1 C= s [41] $end
$var wire 1 D= s [40] $end
$var wire 1 E= s [39] $end
$var wire 1 F= s [38] $end
$var wire 1 G= s [37] $end
$var wire 1 H= s [36] $end
$var wire 1 I= s [35] $end
$var wire 1 J= s [34] $end
$var wire 1 K= s [33] $end
$var wire 1 L= s [32] $end
$var wire 1 M= s [31] $end
$var wire 1 N= s [30] $end
$var wire 1 O= s [29] $end
$var wire 1 P= s [28] $end
$var wire 1 Q= s [27] $end
$var wire 1 R= s [26] $end
$var wire 1 S= s [25] $end
$var wire 1 T= s [24] $end
$var wire 1 U= s [23] $end
$var wire 1 V= s [22] $end
$var wire 1 W= s [21] $end
$var wire 1 X= s [20] $end
$var wire 1 Y= s [19] $end
$var wire 1 Z= s [18] $end
$var wire 1 [= s [17] $end
$var wire 1 \= s [16] $end
$var wire 1 ]= s [15] $end
$var wire 1 ^= s [14] $end
$var wire 1 _= s [13] $end
$var wire 1 `= s [12] $end
$var wire 1 a= s [11] $end
$var wire 1 b= s [10] $end
$var wire 1 c= s [9] $end
$var wire 1 d= s [8] $end
$var wire 1 e= s [7] $end
$var wire 1 f= s [6] $end
$var wire 1 g= s [5] $end
$var wire 1 h= s [4] $end
$var wire 1 i= s [3] $end
$var wire 1 j= s [2] $end
$var wire 1 k= s [1] $end
$var wire 1 l= s [0] $end
$var wire 1 m= ca [42] $end
$var wire 1 n= ca [41] $end
$var wire 1 o= ca [40] $end
$var wire 1 p= ca [39] $end
$var wire 1 q= ca [38] $end
$var wire 1 r= ca [37] $end
$var wire 1 s= ca [36] $end
$var wire 1 t= ca [35] $end
$var wire 1 u= ca [34] $end
$var wire 1 v= ca [33] $end
$var wire 1 w= ca [32] $end
$var wire 1 x= ca [31] $end
$var wire 1 y= ca [30] $end
$var wire 1 z= ca [29] $end
$var wire 1 {= ca [28] $end
$var wire 1 |= ca [27] $end
$var wire 1 }= ca [26] $end
$var wire 1 ~= ca [25] $end
$var wire 1 !> ca [24] $end
$var wire 1 "> ca [23] $end
$var wire 1 #> ca [22] $end
$var wire 1 $> ca [21] $end
$var wire 1 %> ca [20] $end
$var wire 1 &> ca [19] $end
$var wire 1 '> ca [18] $end
$var wire 1 (> ca [17] $end
$var wire 1 )> ca [16] $end
$var wire 1 *> ca [15] $end
$var wire 1 +> ca [14] $end
$var wire 1 ,> ca [13] $end
$var wire 1 -> ca [12] $end
$var wire 1 .> ca [11] $end
$var wire 1 /> ca [10] $end
$var wire 1 0> ca [9] $end
$var wire 1 1> ca [8] $end
$var wire 1 2> ca [7] $end
$var wire 1 3> ca [6] $end
$var wire 1 4> ca [5] $end
$var wire 1 5> ca [4] $end
$var wire 1 6> ca [3] $end
$var wire 1 7> ca [2] $end
$var wire 1 8> ca [1] $end
$var wire 1 9> ca [0] $end
$upscope $end

$scope module l2_2 $end
$var parameter 32 GS size $end
$var wire 1 HS p1 [46] $end
$var wire 1 IS p1 [45] $end
$var wire 1 JS p1 [44] $end
$var wire 1 KS p1 [43] $end
$var wire 1 LS p1 [42] $end
$var wire 1 MS p1 [41] $end
$var wire 1 NS p1 [40] $end
$var wire 1 OS p1 [39] $end
$var wire 1 PS p1 [38] $end
$var wire 1 QS p1 [37] $end
$var wire 1 RS p1 [36] $end
$var wire 1 SS p1 [35] $end
$var wire 1 TS p1 [34] $end
$var wire 1 US p1 [33] $end
$var wire 1 VS p1 [32] $end
$var wire 1 WS p1 [31] $end
$var wire 1 XS p1 [30] $end
$var wire 1 YS p1 [29] $end
$var wire 1 ZS p1 [28] $end
$var wire 1 [S p1 [27] $end
$var wire 1 \S p1 [26] $end
$var wire 1 ]S p1 [25] $end
$var wire 1 ^S p1 [24] $end
$var wire 1 _S p1 [23] $end
$var wire 1 `S p1 [22] $end
$var wire 1 aS p1 [21] $end
$var wire 1 bS p1 [20] $end
$var wire 1 cS p1 [19] $end
$var wire 1 dS p1 [18] $end
$var wire 1 eS p1 [17] $end
$var wire 1 fS p1 [16] $end
$var wire 1 gS p1 [15] $end
$var wire 1 hS p1 [14] $end
$var wire 1 iS p1 [13] $end
$var wire 1 jS p1 [12] $end
$var wire 1 kS p1 [11] $end
$var wire 1 lS p1 [10] $end
$var wire 1 mS p1 [9] $end
$var wire 1 nS p1 [8] $end
$var wire 1 oS p1 [7] $end
$var wire 1 pS p1 [6] $end
$var wire 1 qS p1 [5] $end
$var wire 1 rS p1 [4] $end
$var wire 1 sS p1 [3] $end
$var wire 1 tS p1 [2] $end
$var wire 1 uS p1 [1] $end
$var wire 1 vS p1 [0] $end
$var wire 1 wS p2 [46] $end
$var wire 1 xS p2 [45] $end
$var wire 1 yS p2 [44] $end
$var wire 1 zS p2 [43] $end
$var wire 1 {S p2 [42] $end
$var wire 1 |S p2 [41] $end
$var wire 1 }S p2 [40] $end
$var wire 1 ~S p2 [39] $end
$var wire 1 !T p2 [38] $end
$var wire 1 "T p2 [37] $end
$var wire 1 #T p2 [36] $end
$var wire 1 $T p2 [35] $end
$var wire 1 %T p2 [34] $end
$var wire 1 &T p2 [33] $end
$var wire 1 'T p2 [32] $end
$var wire 1 (T p2 [31] $end
$var wire 1 )T p2 [30] $end
$var wire 1 *T p2 [29] $end
$var wire 1 +T p2 [28] $end
$var wire 1 ,T p2 [27] $end
$var wire 1 -T p2 [26] $end
$var wire 1 .T p2 [25] $end
$var wire 1 /T p2 [24] $end
$var wire 1 0T p2 [23] $end
$var wire 1 1T p2 [22] $end
$var wire 1 2T p2 [21] $end
$var wire 1 3T p2 [20] $end
$var wire 1 4T p2 [19] $end
$var wire 1 5T p2 [18] $end
$var wire 1 6T p2 [17] $end
$var wire 1 7T p2 [16] $end
$var wire 1 8T p2 [15] $end
$var wire 1 9T p2 [14] $end
$var wire 1 :T p2 [13] $end
$var wire 1 ;T p2 [12] $end
$var wire 1 <T p2 [11] $end
$var wire 1 =T p2 [10] $end
$var wire 1 >T p2 [9] $end
$var wire 1 ?T p2 [8] $end
$var wire 1 @T p2 [7] $end
$var wire 1 AT p2 [6] $end
$var wire 1 BT p2 [5] $end
$var wire 1 CT p2 [4] $end
$var wire 1 DT p2 [3] $end
$var wire 1 ET p2 [2] $end
$var wire 1 FT p2 [1] $end
$var wire 1 GT p2 [0] $end
$var wire 1 HT p3 [46] $end
$var wire 1 IT p3 [45] $end
$var wire 1 JT p3 [44] $end
$var wire 1 KT p3 [43] $end
$var wire 1 LT p3 [42] $end
$var wire 1 MT p3 [41] $end
$var wire 1 NT p3 [40] $end
$var wire 1 OT p3 [39] $end
$var wire 1 PT p3 [38] $end
$var wire 1 QT p3 [37] $end
$var wire 1 RT p3 [36] $end
$var wire 1 ST p3 [35] $end
$var wire 1 TT p3 [34] $end
$var wire 1 UT p3 [33] $end
$var wire 1 VT p3 [32] $end
$var wire 1 WT p3 [31] $end
$var wire 1 XT p3 [30] $end
$var wire 1 YT p3 [29] $end
$var wire 1 ZT p3 [28] $end
$var wire 1 [T p3 [27] $end
$var wire 1 \T p3 [26] $end
$var wire 1 ]T p3 [25] $end
$var wire 1 ^T p3 [24] $end
$var wire 1 _T p3 [23] $end
$var wire 1 `T p3 [22] $end
$var wire 1 aT p3 [21] $end
$var wire 1 bT p3 [20] $end
$var wire 1 cT p3 [19] $end
$var wire 1 dT p3 [18] $end
$var wire 1 eT p3 [17] $end
$var wire 1 fT p3 [16] $end
$var wire 1 gT p3 [15] $end
$var wire 1 hT p3 [14] $end
$var wire 1 iT p3 [13] $end
$var wire 1 jT p3 [12] $end
$var wire 1 kT p3 [11] $end
$var wire 1 lT p3 [10] $end
$var wire 1 mT p3 [9] $end
$var wire 1 nT p3 [8] $end
$var wire 1 oT p3 [7] $end
$var wire 1 pT p3 [6] $end
$var wire 1 qT p3 [5] $end
$var wire 1 rT p3 [4] $end
$var wire 1 sT p3 [3] $end
$var wire 1 tT p3 [2] $end
$var wire 1 uT p3 [1] $end
$var wire 1 vT p3 [0] $end
$var wire 1 :> c1 [46] $end
$var wire 1 ;> c1 [45] $end
$var wire 1 <> c1 [44] $end
$var wire 1 => c1 [43] $end
$var wire 1 >> c1 [42] $end
$var wire 1 ?> c1 [41] $end
$var wire 1 @> c1 [40] $end
$var wire 1 A> c1 [39] $end
$var wire 1 B> c1 [38] $end
$var wire 1 C> c1 [37] $end
$var wire 1 D> c1 [36] $end
$var wire 1 E> c1 [35] $end
$var wire 1 F> c1 [34] $end
$var wire 1 G> c1 [33] $end
$var wire 1 H> c1 [32] $end
$var wire 1 I> c1 [31] $end
$var wire 1 J> c1 [30] $end
$var wire 1 K> c1 [29] $end
$var wire 1 L> c1 [28] $end
$var wire 1 M> c1 [27] $end
$var wire 1 N> c1 [26] $end
$var wire 1 O> c1 [25] $end
$var wire 1 P> c1 [24] $end
$var wire 1 Q> c1 [23] $end
$var wire 1 R> c1 [22] $end
$var wire 1 S> c1 [21] $end
$var wire 1 T> c1 [20] $end
$var wire 1 U> c1 [19] $end
$var wire 1 V> c1 [18] $end
$var wire 1 W> c1 [17] $end
$var wire 1 X> c1 [16] $end
$var wire 1 Y> c1 [15] $end
$var wire 1 Z> c1 [14] $end
$var wire 1 [> c1 [13] $end
$var wire 1 \> c1 [12] $end
$var wire 1 ]> c1 [11] $end
$var wire 1 ^> c1 [10] $end
$var wire 1 _> c1 [9] $end
$var wire 1 `> c1 [8] $end
$var wire 1 a> c1 [7] $end
$var wire 1 b> c1 [6] $end
$var wire 1 c> c1 [5] $end
$var wire 1 d> c1 [4] $end
$var wire 1 e> c1 [3] $end
$var wire 1 f> c1 [2] $end
$var wire 1 g> c1 [1] $end
$var wire 1 h> c1 [0] $end
$var wire 1 i> c2 [46] $end
$var wire 1 j> c2 [45] $end
$var wire 1 k> c2 [44] $end
$var wire 1 l> c2 [43] $end
$var wire 1 m> c2 [42] $end
$var wire 1 n> c2 [41] $end
$var wire 1 o> c2 [40] $end
$var wire 1 p> c2 [39] $end
$var wire 1 q> c2 [38] $end
$var wire 1 r> c2 [37] $end
$var wire 1 s> c2 [36] $end
$var wire 1 t> c2 [35] $end
$var wire 1 u> c2 [34] $end
$var wire 1 v> c2 [33] $end
$var wire 1 w> c2 [32] $end
$var wire 1 x> c2 [31] $end
$var wire 1 y> c2 [30] $end
$var wire 1 z> c2 [29] $end
$var wire 1 {> c2 [28] $end
$var wire 1 |> c2 [27] $end
$var wire 1 }> c2 [26] $end
$var wire 1 ~> c2 [25] $end
$var wire 1 !? c2 [24] $end
$var wire 1 "? c2 [23] $end
$var wire 1 #? c2 [22] $end
$var wire 1 $? c2 [21] $end
$var wire 1 %? c2 [20] $end
$var wire 1 &? c2 [19] $end
$var wire 1 '? c2 [18] $end
$var wire 1 (? c2 [17] $end
$var wire 1 )? c2 [16] $end
$var wire 1 *? c2 [15] $end
$var wire 1 +? c2 [14] $end
$var wire 1 ,? c2 [13] $end
$var wire 1 -? c2 [12] $end
$var wire 1 .? c2 [11] $end
$var wire 1 /? c2 [10] $end
$var wire 1 0? c2 [9] $end
$var wire 1 1? c2 [8] $end
$var wire 1 2? c2 [7] $end
$var wire 1 3? c2 [6] $end
$var wire 1 4? c2 [5] $end
$var wire 1 5? c2 [4] $end
$var wire 1 6? c2 [3] $end
$var wire 1 7? c2 [2] $end
$var wire 1 8? c2 [1] $end
$var wire 1 9? c2 [0] $end
$var wire 1 :? c3 [46] $end
$var wire 1 ;? c3 [45] $end
$var wire 1 <? c3 [44] $end
$var wire 1 =? c3 [43] $end
$var wire 1 >? c3 [42] $end
$var wire 1 ?? c3 [41] $end
$var wire 1 @? c3 [40] $end
$var wire 1 A? c3 [39] $end
$var wire 1 B? c3 [38] $end
$var wire 1 C? c3 [37] $end
$var wire 1 D? c3 [36] $end
$var wire 1 E? c3 [35] $end
$var wire 1 F? c3 [34] $end
$var wire 1 G? c3 [33] $end
$var wire 1 H? c3 [32] $end
$var wire 1 I? c3 [31] $end
$var wire 1 J? c3 [30] $end
$var wire 1 K? c3 [29] $end
$var wire 1 L? c3 [28] $end
$var wire 1 M? c3 [27] $end
$var wire 1 N? c3 [26] $end
$var wire 1 O? c3 [25] $end
$var wire 1 P? c3 [24] $end
$var wire 1 Q? c3 [23] $end
$var wire 1 R? c3 [22] $end
$var wire 1 S? c3 [21] $end
$var wire 1 T? c3 [20] $end
$var wire 1 U? c3 [19] $end
$var wire 1 V? c3 [18] $end
$var wire 1 W? c3 [17] $end
$var wire 1 X? c3 [16] $end
$var wire 1 Y? c3 [15] $end
$var wire 1 Z? c3 [14] $end
$var wire 1 [? c3 [13] $end
$var wire 1 \? c3 [12] $end
$var wire 1 ]? c3 [11] $end
$var wire 1 ^? c3 [10] $end
$var wire 1 _? c3 [9] $end
$var wire 1 `? c3 [8] $end
$var wire 1 a? c3 [7] $end
$var wire 1 b? c3 [6] $end
$var wire 1 c? c3 [5] $end
$var wire 1 d? c3 [4] $end
$var wire 1 e? c3 [3] $end
$var wire 1 f? c3 [2] $end
$var wire 1 g? c3 [1] $end
$var wire 1 h? c3 [0] $end
$var wire 1 i? c4 [46] $end
$var wire 1 j? c4 [45] $end
$var wire 1 k? c4 [44] $end
$var wire 1 l? c4 [43] $end
$var wire 1 m? c4 [42] $end
$var wire 1 n? c4 [41] $end
$var wire 1 o? c4 [40] $end
$var wire 1 p? c4 [39] $end
$var wire 1 q? c4 [38] $end
$var wire 1 r? c4 [37] $end
$var wire 1 s? c4 [36] $end
$var wire 1 t? c4 [35] $end
$var wire 1 u? c4 [34] $end
$var wire 1 v? c4 [33] $end
$var wire 1 w? c4 [32] $end
$var wire 1 x? c4 [31] $end
$var wire 1 y? c4 [30] $end
$var wire 1 z? c4 [29] $end
$var wire 1 {? c4 [28] $end
$var wire 1 |? c4 [27] $end
$var wire 1 }? c4 [26] $end
$var wire 1 ~? c4 [25] $end
$var wire 1 !@ c4 [24] $end
$var wire 1 "@ c4 [23] $end
$var wire 1 #@ c4 [22] $end
$var wire 1 $@ c4 [21] $end
$var wire 1 %@ c4 [20] $end
$var wire 1 &@ c4 [19] $end
$var wire 1 '@ c4 [18] $end
$var wire 1 (@ c4 [17] $end
$var wire 1 )@ c4 [16] $end
$var wire 1 *@ c4 [15] $end
$var wire 1 +@ c4 [14] $end
$var wire 1 ,@ c4 [13] $end
$var wire 1 -@ c4 [12] $end
$var wire 1 .@ c4 [11] $end
$var wire 1 /@ c4 [10] $end
$var wire 1 0@ c4 [9] $end
$var wire 1 1@ c4 [8] $end
$var wire 1 2@ c4 [7] $end
$var wire 1 3@ c4 [6] $end
$var wire 1 4@ c4 [5] $end
$var wire 1 5@ c4 [4] $end
$var wire 1 6@ c4 [3] $end
$var wire 1 7@ c4 [2] $end
$var wire 1 8@ c4 [1] $end
$var wire 1 9@ c4 [0] $end
$var wire 1 :@ cin [46] $end
$var wire 1 ;@ cin [45] $end
$var wire 1 <@ cin [44] $end
$var wire 1 =@ cin [43] $end
$var wire 1 >@ cin [42] $end
$var wire 1 ?@ cin [41] $end
$var wire 1 @@ cin [40] $end
$var wire 1 A@ cin [39] $end
$var wire 1 B@ cin [38] $end
$var wire 1 C@ cin [37] $end
$var wire 1 D@ cin [36] $end
$var wire 1 E@ cin [35] $end
$var wire 1 F@ cin [34] $end
$var wire 1 G@ cin [33] $end
$var wire 1 H@ cin [32] $end
$var wire 1 I@ cin [31] $end
$var wire 1 J@ cin [30] $end
$var wire 1 K@ cin [29] $end
$var wire 1 L@ cin [28] $end
$var wire 1 M@ cin [27] $end
$var wire 1 N@ cin [26] $end
$var wire 1 O@ cin [25] $end
$var wire 1 P@ cin [24] $end
$var wire 1 Q@ cin [23] $end
$var wire 1 R@ cin [22] $end
$var wire 1 S@ cin [21] $end
$var wire 1 T@ cin [20] $end
$var wire 1 U@ cin [19] $end
$var wire 1 V@ cin [18] $end
$var wire 1 W@ cin [17] $end
$var wire 1 X@ cin [16] $end
$var wire 1 Y@ cin [15] $end
$var wire 1 Z@ cin [14] $end
$var wire 1 [@ cin [13] $end
$var wire 1 \@ cin [12] $end
$var wire 1 ]@ cin [11] $end
$var wire 1 ^@ cin [10] $end
$var wire 1 _@ cin [9] $end
$var wire 1 `@ cin [8] $end
$var wire 1 a@ cin [7] $end
$var wire 1 b@ cin [6] $end
$var wire 1 c@ cin [5] $end
$var wire 1 d@ cin [4] $end
$var wire 1 e@ cin [3] $end
$var wire 1 f@ cin [2] $end
$var wire 1 g@ cin [1] $end
$var wire 1 h@ cin [0] $end
$var wire 1 i@ cout [46] $end
$var wire 1 j@ cout [45] $end
$var wire 1 k@ cout [44] $end
$var wire 1 l@ cout [43] $end
$var wire 1 m@ cout [42] $end
$var wire 1 n@ cout [41] $end
$var wire 1 o@ cout [40] $end
$var wire 1 p@ cout [39] $end
$var wire 1 q@ cout [38] $end
$var wire 1 r@ cout [37] $end
$var wire 1 s@ cout [36] $end
$var wire 1 t@ cout [35] $end
$var wire 1 u@ cout [34] $end
$var wire 1 v@ cout [33] $end
$var wire 1 w@ cout [32] $end
$var wire 1 x@ cout [31] $end
$var wire 1 y@ cout [30] $end
$var wire 1 z@ cout [29] $end
$var wire 1 {@ cout [28] $end
$var wire 1 |@ cout [27] $end
$var wire 1 }@ cout [26] $end
$var wire 1 ~@ cout [25] $end
$var wire 1 !A cout [24] $end
$var wire 1 "A cout [23] $end
$var wire 1 #A cout [22] $end
$var wire 1 $A cout [21] $end
$var wire 1 %A cout [20] $end
$var wire 1 &A cout [19] $end
$var wire 1 'A cout [18] $end
$var wire 1 (A cout [17] $end
$var wire 1 )A cout [16] $end
$var wire 1 *A cout [15] $end
$var wire 1 +A cout [14] $end
$var wire 1 ,A cout [13] $end
$var wire 1 -A cout [12] $end
$var wire 1 .A cout [11] $end
$var wire 1 /A cout [10] $end
$var wire 1 0A cout [9] $end
$var wire 1 1A cout [8] $end
$var wire 1 2A cout [7] $end
$var wire 1 3A cout [6] $end
$var wire 1 4A cout [5] $end
$var wire 1 5A cout [4] $end
$var wire 1 6A cout [3] $end
$var wire 1 7A cout [2] $end
$var wire 1 8A cout [1] $end
$var wire 1 9A cout [0] $end
$var wire 1 :A s [46] $end
$var wire 1 ;A s [45] $end
$var wire 1 <A s [44] $end
$var wire 1 =A s [43] $end
$var wire 1 >A s [42] $end
$var wire 1 ?A s [41] $end
$var wire 1 @A s [40] $end
$var wire 1 AA s [39] $end
$var wire 1 BA s [38] $end
$var wire 1 CA s [37] $end
$var wire 1 DA s [36] $end
$var wire 1 EA s [35] $end
$var wire 1 FA s [34] $end
$var wire 1 GA s [33] $end
$var wire 1 HA s [32] $end
$var wire 1 IA s [31] $end
$var wire 1 JA s [30] $end
$var wire 1 KA s [29] $end
$var wire 1 LA s [28] $end
$var wire 1 MA s [27] $end
$var wire 1 NA s [26] $end
$var wire 1 OA s [25] $end
$var wire 1 PA s [24] $end
$var wire 1 QA s [23] $end
$var wire 1 RA s [22] $end
$var wire 1 SA s [21] $end
$var wire 1 TA s [20] $end
$var wire 1 UA s [19] $end
$var wire 1 VA s [18] $end
$var wire 1 WA s [17] $end
$var wire 1 XA s [16] $end
$var wire 1 YA s [15] $end
$var wire 1 ZA s [14] $end
$var wire 1 [A s [13] $end
$var wire 1 \A s [12] $end
$var wire 1 ]A s [11] $end
$var wire 1 ^A s [10] $end
$var wire 1 _A s [9] $end
$var wire 1 `A s [8] $end
$var wire 1 aA s [7] $end
$var wire 1 bA s [6] $end
$var wire 1 cA s [5] $end
$var wire 1 dA s [4] $end
$var wire 1 eA s [3] $end
$var wire 1 fA s [2] $end
$var wire 1 gA s [1] $end
$var wire 1 hA s [0] $end
$var wire 1 iA ca [46] $end
$var wire 1 jA ca [45] $end
$var wire 1 kA ca [44] $end
$var wire 1 lA ca [43] $end
$var wire 1 mA ca [42] $end
$var wire 1 nA ca [41] $end
$var wire 1 oA ca [40] $end
$var wire 1 pA ca [39] $end
$var wire 1 qA ca [38] $end
$var wire 1 rA ca [37] $end
$var wire 1 sA ca [36] $end
$var wire 1 tA ca [35] $end
$var wire 1 uA ca [34] $end
$var wire 1 vA ca [33] $end
$var wire 1 wA ca [32] $end
$var wire 1 xA ca [31] $end
$var wire 1 yA ca [30] $end
$var wire 1 zA ca [29] $end
$var wire 1 {A ca [28] $end
$var wire 1 |A ca [27] $end
$var wire 1 }A ca [26] $end
$var wire 1 ~A ca [25] $end
$var wire 1 !B ca [24] $end
$var wire 1 "B ca [23] $end
$var wire 1 #B ca [22] $end
$var wire 1 $B ca [21] $end
$var wire 1 %B ca [20] $end
$var wire 1 &B ca [19] $end
$var wire 1 'B ca [18] $end
$var wire 1 (B ca [17] $end
$var wire 1 )B ca [16] $end
$var wire 1 *B ca [15] $end
$var wire 1 +B ca [14] $end
$var wire 1 ,B ca [13] $end
$var wire 1 -B ca [12] $end
$var wire 1 .B ca [11] $end
$var wire 1 /B ca [10] $end
$var wire 1 0B ca [9] $end
$var wire 1 1B ca [8] $end
$var wire 1 2B ca [7] $end
$var wire 1 3B ca [6] $end
$var wire 1 4B ca [5] $end
$var wire 1 5B ca [4] $end
$var wire 1 6B ca [3] $end
$var wire 1 7B ca [2] $end
$var wire 1 8B ca [1] $end
$var wire 1 9B ca [0] $end
$upscope $end

$scope module l2_3 $end
$var parameter 32 wT size $end
$var wire 1 xT p1 [43] $end
$var wire 1 yT p1 [42] $end
$var wire 1 zT p1 [41] $end
$var wire 1 {T p1 [40] $end
$var wire 1 |T p1 [39] $end
$var wire 1 }T p1 [38] $end
$var wire 1 ~T p1 [37] $end
$var wire 1 !U p1 [36] $end
$var wire 1 "U p1 [35] $end
$var wire 1 #U p1 [34] $end
$var wire 1 $U p1 [33] $end
$var wire 1 %U p1 [32] $end
$var wire 1 &U p1 [31] $end
$var wire 1 'U p1 [30] $end
$var wire 1 (U p1 [29] $end
$var wire 1 )U p1 [28] $end
$var wire 1 *U p1 [27] $end
$var wire 1 +U p1 [26] $end
$var wire 1 ,U p1 [25] $end
$var wire 1 -U p1 [24] $end
$var wire 1 .U p1 [23] $end
$var wire 1 /U p1 [22] $end
$var wire 1 0U p1 [21] $end
$var wire 1 1U p1 [20] $end
$var wire 1 2U p1 [19] $end
$var wire 1 3U p1 [18] $end
$var wire 1 4U p1 [17] $end
$var wire 1 5U p1 [16] $end
$var wire 1 6U p1 [15] $end
$var wire 1 7U p1 [14] $end
$var wire 1 8U p1 [13] $end
$var wire 1 9U p1 [12] $end
$var wire 1 :U p1 [11] $end
$var wire 1 ;U p1 [10] $end
$var wire 1 <U p1 [9] $end
$var wire 1 =U p1 [8] $end
$var wire 1 >U p1 [7] $end
$var wire 1 ?U p1 [6] $end
$var wire 1 @U p1 [5] $end
$var wire 1 AU p1 [4] $end
$var wire 1 BU p1 [3] $end
$var wire 1 CU p1 [2] $end
$var wire 1 DU p1 [1] $end
$var wire 1 EU p1 [0] $end
$var wire 1 FU p2 [43] $end
$var wire 1 GU p2 [42] $end
$var wire 1 HU p2 [41] $end
$var wire 1 IU p2 [40] $end
$var wire 1 JU p2 [39] $end
$var wire 1 KU p2 [38] $end
$var wire 1 LU p2 [37] $end
$var wire 1 MU p2 [36] $end
$var wire 1 NU p2 [35] $end
$var wire 1 OU p2 [34] $end
$var wire 1 PU p2 [33] $end
$var wire 1 QU p2 [32] $end
$var wire 1 RU p2 [31] $end
$var wire 1 SU p2 [30] $end
$var wire 1 TU p2 [29] $end
$var wire 1 UU p2 [28] $end
$var wire 1 VU p2 [27] $end
$var wire 1 WU p2 [26] $end
$var wire 1 XU p2 [25] $end
$var wire 1 YU p2 [24] $end
$var wire 1 ZU p2 [23] $end
$var wire 1 [U p2 [22] $end
$var wire 1 \U p2 [21] $end
$var wire 1 ]U p2 [20] $end
$var wire 1 ^U p2 [19] $end
$var wire 1 _U p2 [18] $end
$var wire 1 `U p2 [17] $end
$var wire 1 aU p2 [16] $end
$var wire 1 bU p2 [15] $end
$var wire 1 cU p2 [14] $end
$var wire 1 dU p2 [13] $end
$var wire 1 eU p2 [12] $end
$var wire 1 fU p2 [11] $end
$var wire 1 gU p2 [10] $end
$var wire 1 hU p2 [9] $end
$var wire 1 iU p2 [8] $end
$var wire 1 jU p2 [7] $end
$var wire 1 kU p2 [6] $end
$var wire 1 lU p2 [5] $end
$var wire 1 mU p2 [4] $end
$var wire 1 nU p2 [3] $end
$var wire 1 oU p2 [2] $end
$var wire 1 pU p2 [1] $end
$var wire 1 qU p2 [0] $end
$var wire 1 rU p3 [43] $end
$var wire 1 sU p3 [42] $end
$var wire 1 tU p3 [41] $end
$var wire 1 uU p3 [40] $end
$var wire 1 vU p3 [39] $end
$var wire 1 wU p3 [38] $end
$var wire 1 xU p3 [37] $end
$var wire 1 yU p3 [36] $end
$var wire 1 zU p3 [35] $end
$var wire 1 {U p3 [34] $end
$var wire 1 |U p3 [33] $end
$var wire 1 }U p3 [32] $end
$var wire 1 ~U p3 [31] $end
$var wire 1 !V p3 [30] $end
$var wire 1 "V p3 [29] $end
$var wire 1 #V p3 [28] $end
$var wire 1 $V p3 [27] $end
$var wire 1 %V p3 [26] $end
$var wire 1 &V p3 [25] $end
$var wire 1 'V p3 [24] $end
$var wire 1 (V p3 [23] $end
$var wire 1 )V p3 [22] $end
$var wire 1 *V p3 [21] $end
$var wire 1 +V p3 [20] $end
$var wire 1 ,V p3 [19] $end
$var wire 1 -V p3 [18] $end
$var wire 1 .V p3 [17] $end
$var wire 1 /V p3 [16] $end
$var wire 1 0V p3 [15] $end
$var wire 1 1V p3 [14] $end
$var wire 1 2V p3 [13] $end
$var wire 1 3V p3 [12] $end
$var wire 1 4V p3 [11] $end
$var wire 1 5V p3 [10] $end
$var wire 1 6V p3 [9] $end
$var wire 1 7V p3 [8] $end
$var wire 1 8V p3 [7] $end
$var wire 1 9V p3 [6] $end
$var wire 1 :V p3 [5] $end
$var wire 1 ;V p3 [4] $end
$var wire 1 <V p3 [3] $end
$var wire 1 =V p3 [2] $end
$var wire 1 >V p3 [1] $end
$var wire 1 ?V p3 [0] $end
$var wire 1 :B c1 [43] $end
$var wire 1 ;B c1 [42] $end
$var wire 1 <B c1 [41] $end
$var wire 1 =B c1 [40] $end
$var wire 1 >B c1 [39] $end
$var wire 1 ?B c1 [38] $end
$var wire 1 @B c1 [37] $end
$var wire 1 AB c1 [36] $end
$var wire 1 BB c1 [35] $end
$var wire 1 CB c1 [34] $end
$var wire 1 DB c1 [33] $end
$var wire 1 EB c1 [32] $end
$var wire 1 FB c1 [31] $end
$var wire 1 GB c1 [30] $end
$var wire 1 HB c1 [29] $end
$var wire 1 IB c1 [28] $end
$var wire 1 JB c1 [27] $end
$var wire 1 KB c1 [26] $end
$var wire 1 LB c1 [25] $end
$var wire 1 MB c1 [24] $end
$var wire 1 NB c1 [23] $end
$var wire 1 OB c1 [22] $end
$var wire 1 PB c1 [21] $end
$var wire 1 QB c1 [20] $end
$var wire 1 RB c1 [19] $end
$var wire 1 SB c1 [18] $end
$var wire 1 TB c1 [17] $end
$var wire 1 UB c1 [16] $end
$var wire 1 VB c1 [15] $end
$var wire 1 WB c1 [14] $end
$var wire 1 XB c1 [13] $end
$var wire 1 YB c1 [12] $end
$var wire 1 ZB c1 [11] $end
$var wire 1 [B c1 [10] $end
$var wire 1 \B c1 [9] $end
$var wire 1 ]B c1 [8] $end
$var wire 1 ^B c1 [7] $end
$var wire 1 _B c1 [6] $end
$var wire 1 `B c1 [5] $end
$var wire 1 aB c1 [4] $end
$var wire 1 bB c1 [3] $end
$var wire 1 cB c1 [2] $end
$var wire 1 dB c1 [1] $end
$var wire 1 eB c1 [0] $end
$var wire 1 fB c2 [43] $end
$var wire 1 gB c2 [42] $end
$var wire 1 hB c2 [41] $end
$var wire 1 iB c2 [40] $end
$var wire 1 jB c2 [39] $end
$var wire 1 kB c2 [38] $end
$var wire 1 lB c2 [37] $end
$var wire 1 mB c2 [36] $end
$var wire 1 nB c2 [35] $end
$var wire 1 oB c2 [34] $end
$var wire 1 pB c2 [33] $end
$var wire 1 qB c2 [32] $end
$var wire 1 rB c2 [31] $end
$var wire 1 sB c2 [30] $end
$var wire 1 tB c2 [29] $end
$var wire 1 uB c2 [28] $end
$var wire 1 vB c2 [27] $end
$var wire 1 wB c2 [26] $end
$var wire 1 xB c2 [25] $end
$var wire 1 yB c2 [24] $end
$var wire 1 zB c2 [23] $end
$var wire 1 {B c2 [22] $end
$var wire 1 |B c2 [21] $end
$var wire 1 }B c2 [20] $end
$var wire 1 ~B c2 [19] $end
$var wire 1 !C c2 [18] $end
$var wire 1 "C c2 [17] $end
$var wire 1 #C c2 [16] $end
$var wire 1 $C c2 [15] $end
$var wire 1 %C c2 [14] $end
$var wire 1 &C c2 [13] $end
$var wire 1 'C c2 [12] $end
$var wire 1 (C c2 [11] $end
$var wire 1 )C c2 [10] $end
$var wire 1 *C c2 [9] $end
$var wire 1 +C c2 [8] $end
$var wire 1 ,C c2 [7] $end
$var wire 1 -C c2 [6] $end
$var wire 1 .C c2 [5] $end
$var wire 1 /C c2 [4] $end
$var wire 1 0C c2 [3] $end
$var wire 1 1C c2 [2] $end
$var wire 1 2C c2 [1] $end
$var wire 1 3C c2 [0] $end
$var wire 1 4C c3 [43] $end
$var wire 1 5C c3 [42] $end
$var wire 1 6C c3 [41] $end
$var wire 1 7C c3 [40] $end
$var wire 1 8C c3 [39] $end
$var wire 1 9C c3 [38] $end
$var wire 1 :C c3 [37] $end
$var wire 1 ;C c3 [36] $end
$var wire 1 <C c3 [35] $end
$var wire 1 =C c3 [34] $end
$var wire 1 >C c3 [33] $end
$var wire 1 ?C c3 [32] $end
$var wire 1 @C c3 [31] $end
$var wire 1 AC c3 [30] $end
$var wire 1 BC c3 [29] $end
$var wire 1 CC c3 [28] $end
$var wire 1 DC c3 [27] $end
$var wire 1 EC c3 [26] $end
$var wire 1 FC c3 [25] $end
$var wire 1 GC c3 [24] $end
$var wire 1 HC c3 [23] $end
$var wire 1 IC c3 [22] $end
$var wire 1 JC c3 [21] $end
$var wire 1 KC c3 [20] $end
$var wire 1 LC c3 [19] $end
$var wire 1 MC c3 [18] $end
$var wire 1 NC c3 [17] $end
$var wire 1 OC c3 [16] $end
$var wire 1 PC c3 [15] $end
$var wire 1 QC c3 [14] $end
$var wire 1 RC c3 [13] $end
$var wire 1 SC c3 [12] $end
$var wire 1 TC c3 [11] $end
$var wire 1 UC c3 [10] $end
$var wire 1 VC c3 [9] $end
$var wire 1 WC c3 [8] $end
$var wire 1 XC c3 [7] $end
$var wire 1 YC c3 [6] $end
$var wire 1 ZC c3 [5] $end
$var wire 1 [C c3 [4] $end
$var wire 1 \C c3 [3] $end
$var wire 1 ]C c3 [2] $end
$var wire 1 ^C c3 [1] $end
$var wire 1 _C c3 [0] $end
$var wire 1 `C c4 [43] $end
$var wire 1 aC c4 [42] $end
$var wire 1 bC c4 [41] $end
$var wire 1 cC c4 [40] $end
$var wire 1 dC c4 [39] $end
$var wire 1 eC c4 [38] $end
$var wire 1 fC c4 [37] $end
$var wire 1 gC c4 [36] $end
$var wire 1 hC c4 [35] $end
$var wire 1 iC c4 [34] $end
$var wire 1 jC c4 [33] $end
$var wire 1 kC c4 [32] $end
$var wire 1 lC c4 [31] $end
$var wire 1 mC c4 [30] $end
$var wire 1 nC c4 [29] $end
$var wire 1 oC c4 [28] $end
$var wire 1 pC c4 [27] $end
$var wire 1 qC c4 [26] $end
$var wire 1 rC c4 [25] $end
$var wire 1 sC c4 [24] $end
$var wire 1 tC c4 [23] $end
$var wire 1 uC c4 [22] $end
$var wire 1 vC c4 [21] $end
$var wire 1 wC c4 [20] $end
$var wire 1 xC c4 [19] $end
$var wire 1 yC c4 [18] $end
$var wire 1 zC c4 [17] $end
$var wire 1 {C c4 [16] $end
$var wire 1 |C c4 [15] $end
$var wire 1 }C c4 [14] $end
$var wire 1 ~C c4 [13] $end
$var wire 1 !D c4 [12] $end
$var wire 1 "D c4 [11] $end
$var wire 1 #D c4 [10] $end
$var wire 1 $D c4 [9] $end
$var wire 1 %D c4 [8] $end
$var wire 1 &D c4 [7] $end
$var wire 1 'D c4 [6] $end
$var wire 1 (D c4 [5] $end
$var wire 1 )D c4 [4] $end
$var wire 1 *D c4 [3] $end
$var wire 1 +D c4 [2] $end
$var wire 1 ,D c4 [1] $end
$var wire 1 -D c4 [0] $end
$var wire 1 .D cin [43] $end
$var wire 1 /D cin [42] $end
$var wire 1 0D cin [41] $end
$var wire 1 1D cin [40] $end
$var wire 1 2D cin [39] $end
$var wire 1 3D cin [38] $end
$var wire 1 4D cin [37] $end
$var wire 1 5D cin [36] $end
$var wire 1 6D cin [35] $end
$var wire 1 7D cin [34] $end
$var wire 1 8D cin [33] $end
$var wire 1 9D cin [32] $end
$var wire 1 :D cin [31] $end
$var wire 1 ;D cin [30] $end
$var wire 1 <D cin [29] $end
$var wire 1 =D cin [28] $end
$var wire 1 >D cin [27] $end
$var wire 1 ?D cin [26] $end
$var wire 1 @D cin [25] $end
$var wire 1 AD cin [24] $end
$var wire 1 BD cin [23] $end
$var wire 1 CD cin [22] $end
$var wire 1 DD cin [21] $end
$var wire 1 ED cin [20] $end
$var wire 1 FD cin [19] $end
$var wire 1 GD cin [18] $end
$var wire 1 HD cin [17] $end
$var wire 1 ID cin [16] $end
$var wire 1 JD cin [15] $end
$var wire 1 KD cin [14] $end
$var wire 1 LD cin [13] $end
$var wire 1 MD cin [12] $end
$var wire 1 ND cin [11] $end
$var wire 1 OD cin [10] $end
$var wire 1 PD cin [9] $end
$var wire 1 QD cin [8] $end
$var wire 1 RD cin [7] $end
$var wire 1 SD cin [6] $end
$var wire 1 TD cin [5] $end
$var wire 1 UD cin [4] $end
$var wire 1 VD cin [3] $end
$var wire 1 WD cin [2] $end
$var wire 1 XD cin [1] $end
$var wire 1 YD cin [0] $end
$var wire 1 ZD cout [43] $end
$var wire 1 [D cout [42] $end
$var wire 1 \D cout [41] $end
$var wire 1 ]D cout [40] $end
$var wire 1 ^D cout [39] $end
$var wire 1 _D cout [38] $end
$var wire 1 `D cout [37] $end
$var wire 1 aD cout [36] $end
$var wire 1 bD cout [35] $end
$var wire 1 cD cout [34] $end
$var wire 1 dD cout [33] $end
$var wire 1 eD cout [32] $end
$var wire 1 fD cout [31] $end
$var wire 1 gD cout [30] $end
$var wire 1 hD cout [29] $end
$var wire 1 iD cout [28] $end
$var wire 1 jD cout [27] $end
$var wire 1 kD cout [26] $end
$var wire 1 lD cout [25] $end
$var wire 1 mD cout [24] $end
$var wire 1 nD cout [23] $end
$var wire 1 oD cout [22] $end
$var wire 1 pD cout [21] $end
$var wire 1 qD cout [20] $end
$var wire 1 rD cout [19] $end
$var wire 1 sD cout [18] $end
$var wire 1 tD cout [17] $end
$var wire 1 uD cout [16] $end
$var wire 1 vD cout [15] $end
$var wire 1 wD cout [14] $end
$var wire 1 xD cout [13] $end
$var wire 1 yD cout [12] $end
$var wire 1 zD cout [11] $end
$var wire 1 {D cout [10] $end
$var wire 1 |D cout [9] $end
$var wire 1 }D cout [8] $end
$var wire 1 ~D cout [7] $end
$var wire 1 !E cout [6] $end
$var wire 1 "E cout [5] $end
$var wire 1 #E cout [4] $end
$var wire 1 $E cout [3] $end
$var wire 1 %E cout [2] $end
$var wire 1 &E cout [1] $end
$var wire 1 'E cout [0] $end
$var wire 1 (E s [43] $end
$var wire 1 )E s [42] $end
$var wire 1 *E s [41] $end
$var wire 1 +E s [40] $end
$var wire 1 ,E s [39] $end
$var wire 1 -E s [38] $end
$var wire 1 .E s [37] $end
$var wire 1 /E s [36] $end
$var wire 1 0E s [35] $end
$var wire 1 1E s [34] $end
$var wire 1 2E s [33] $end
$var wire 1 3E s [32] $end
$var wire 1 4E s [31] $end
$var wire 1 5E s [30] $end
$var wire 1 6E s [29] $end
$var wire 1 7E s [28] $end
$var wire 1 8E s [27] $end
$var wire 1 9E s [26] $end
$var wire 1 :E s [25] $end
$var wire 1 ;E s [24] $end
$var wire 1 <E s [23] $end
$var wire 1 =E s [22] $end
$var wire 1 >E s [21] $end
$var wire 1 ?E s [20] $end
$var wire 1 @E s [19] $end
$var wire 1 AE s [18] $end
$var wire 1 BE s [17] $end
$var wire 1 CE s [16] $end
$var wire 1 DE s [15] $end
$var wire 1 EE s [14] $end
$var wire 1 FE s [13] $end
$var wire 1 GE s [12] $end
$var wire 1 HE s [11] $end
$var wire 1 IE s [10] $end
$var wire 1 JE s [9] $end
$var wire 1 KE s [8] $end
$var wire 1 LE s [7] $end
$var wire 1 ME s [6] $end
$var wire 1 NE s [5] $end
$var wire 1 OE s [4] $end
$var wire 1 PE s [3] $end
$var wire 1 QE s [2] $end
$var wire 1 RE s [1] $end
$var wire 1 SE s [0] $end
$var wire 1 TE ca [43] $end
$var wire 1 UE ca [42] $end
$var wire 1 VE ca [41] $end
$var wire 1 WE ca [40] $end
$var wire 1 XE ca [39] $end
$var wire 1 YE ca [38] $end
$var wire 1 ZE ca [37] $end
$var wire 1 [E ca [36] $end
$var wire 1 \E ca [35] $end
$var wire 1 ]E ca [34] $end
$var wire 1 ^E ca [33] $end
$var wire 1 _E ca [32] $end
$var wire 1 `E ca [31] $end
$var wire 1 aE ca [30] $end
$var wire 1 bE ca [29] $end
$var wire 1 cE ca [28] $end
$var wire 1 dE ca [27] $end
$var wire 1 eE ca [26] $end
$var wire 1 fE ca [25] $end
$var wire 1 gE ca [24] $end
$var wire 1 hE ca [23] $end
$var wire 1 iE ca [22] $end
$var wire 1 jE ca [21] $end
$var wire 1 kE ca [20] $end
$var wire 1 lE ca [19] $end
$var wire 1 mE ca [18] $end
$var wire 1 nE ca [17] $end
$var wire 1 oE ca [16] $end
$var wire 1 pE ca [15] $end
$var wire 1 qE ca [14] $end
$var wire 1 rE ca [13] $end
$var wire 1 sE ca [12] $end
$var wire 1 tE ca [11] $end
$var wire 1 uE ca [10] $end
$var wire 1 vE ca [9] $end
$var wire 1 wE ca [8] $end
$var wire 1 xE ca [7] $end
$var wire 1 yE ca [6] $end
$var wire 1 zE ca [5] $end
$var wire 1 {E ca [4] $end
$var wire 1 |E ca [3] $end
$var wire 1 }E ca [2] $end
$var wire 1 ~E ca [1] $end
$var wire 1 !F ca [0] $end
$upscope $end

$scope module l3_1 $end
$var parameter 32 @V size $end
$var wire 1 (F c0 [54] $end
$var wire 1 )F c0 [53] $end
$var wire 1 *F c0 [52] $end
$var wire 1 +F c0 [51] $end
$var wire 1 ,F c0 [50] $end
$var wire 1 -F c0 [49] $end
$var wire 1 .F c0 [48] $end
$var wire 1 /F c0 [47] $end
$var wire 1 0F c0 [46] $end
$var wire 1 1F c0 [45] $end
$var wire 1 2F c0 [44] $end
$var wire 1 3F c0 [43] $end
$var wire 1 4F c0 [42] $end
$var wire 1 5F c0 [41] $end
$var wire 1 6F c0 [40] $end
$var wire 1 7F c0 [39] $end
$var wire 1 8F c0 [38] $end
$var wire 1 9F c0 [37] $end
$var wire 1 :F c0 [36] $end
$var wire 1 ;F c0 [35] $end
$var wire 1 <F c0 [34] $end
$var wire 1 =F c0 [33] $end
$var wire 1 >F c0 [32] $end
$var wire 1 ?F c0 [31] $end
$var wire 1 @F c0 [30] $end
$var wire 1 AF c0 [29] $end
$var wire 1 BF c0 [28] $end
$var wire 1 CF c0 [27] $end
$var wire 1 DF c0 [26] $end
$var wire 1 EF c0 [25] $end
$var wire 1 FF c0 [24] $end
$var wire 1 GF c0 [23] $end
$var wire 1 HF c0 [22] $end
$var wire 1 IF c0 [21] $end
$var wire 1 JF c0 [20] $end
$var wire 1 KF c0 [19] $end
$var wire 1 LF c0 [18] $end
$var wire 1 MF c0 [17] $end
$var wire 1 NF c0 [16] $end
$var wire 1 OF c0 [15] $end
$var wire 1 PF c0 [14] $end
$var wire 1 QF c0 [13] $end
$var wire 1 RF c0 [12] $end
$var wire 1 SF c0 [11] $end
$var wire 1 TF c0 [10] $end
$var wire 1 UF c0 [9] $end
$var wire 1 VF c0 [8] $end
$var wire 1 WF c0 [7] $end
$var wire 1 XF c0 [6] $end
$var wire 1 YF c0 [5] $end
$var wire 1 ZF c0 [4] $end
$var wire 1 [F c0 [3] $end
$var wire 1 \F c0 [2] $end
$var wire 1 ]F c0 [1] $end
$var wire 1 ^F c0 [0] $end
$var wire 1 _F c1 [54] $end
$var wire 1 `F c1 [53] $end
$var wire 1 aF c1 [52] $end
$var wire 1 bF c1 [51] $end
$var wire 1 cF c1 [50] $end
$var wire 1 dF c1 [49] $end
$var wire 1 eF c1 [48] $end
$var wire 1 fF c1 [47] $end
$var wire 1 gF c1 [46] $end
$var wire 1 hF c1 [45] $end
$var wire 1 iF c1 [44] $end
$var wire 1 jF c1 [43] $end
$var wire 1 kF c1 [42] $end
$var wire 1 lF c1 [41] $end
$var wire 1 mF c1 [40] $end
$var wire 1 nF c1 [39] $end
$var wire 1 oF c1 [38] $end
$var wire 1 pF c1 [37] $end
$var wire 1 qF c1 [36] $end
$var wire 1 rF c1 [35] $end
$var wire 1 sF c1 [34] $end
$var wire 1 tF c1 [33] $end
$var wire 1 uF c1 [32] $end
$var wire 1 vF c1 [31] $end
$var wire 1 wF c1 [30] $end
$var wire 1 xF c1 [29] $end
$var wire 1 yF c1 [28] $end
$var wire 1 zF c1 [27] $end
$var wire 1 {F c1 [26] $end
$var wire 1 |F c1 [25] $end
$var wire 1 }F c1 [24] $end
$var wire 1 ~F c1 [23] $end
$var wire 1 !G c1 [22] $end
$var wire 1 "G c1 [21] $end
$var wire 1 #G c1 [20] $end
$var wire 1 $G c1 [19] $end
$var wire 1 %G c1 [18] $end
$var wire 1 &G c1 [17] $end
$var wire 1 'G c1 [16] $end
$var wire 1 (G c1 [15] $end
$var wire 1 )G c1 [14] $end
$var wire 1 *G c1 [13] $end
$var wire 1 +G c1 [12] $end
$var wire 1 ,G c1 [11] $end
$var wire 1 -G c1 [10] $end
$var wire 1 .G c1 [9] $end
$var wire 1 /G c1 [8] $end
$var wire 1 0G c1 [7] $end
$var wire 1 1G c1 [6] $end
$var wire 1 2G c1 [5] $end
$var wire 1 3G c1 [4] $end
$var wire 1 4G c1 [3] $end
$var wire 1 5G c1 [2] $end
$var wire 1 6G c1 [1] $end
$var wire 1 7G c1 [0] $end
$var wire 1 8G c2 [54] $end
$var wire 1 9G c2 [53] $end
$var wire 1 :G c2 [52] $end
$var wire 1 ;G c2 [51] $end
$var wire 1 <G c2 [50] $end
$var wire 1 =G c2 [49] $end
$var wire 1 >G c2 [48] $end
$var wire 1 ?G c2 [47] $end
$var wire 1 @G c2 [46] $end
$var wire 1 AG c2 [45] $end
$var wire 1 BG c2 [44] $end
$var wire 1 CG c2 [43] $end
$var wire 1 DG c2 [42] $end
$var wire 1 EG c2 [41] $end
$var wire 1 FG c2 [40] $end
$var wire 1 GG c2 [39] $end
$var wire 1 HG c2 [38] $end
$var wire 1 IG c2 [37] $end
$var wire 1 JG c2 [36] $end
$var wire 1 KG c2 [35] $end
$var wire 1 LG c2 [34] $end
$var wire 1 MG c2 [33] $end
$var wire 1 NG c2 [32] $end
$var wire 1 OG c2 [31] $end
$var wire 1 PG c2 [30] $end
$var wire 1 QG c2 [29] $end
$var wire 1 RG c2 [28] $end
$var wire 1 SG c2 [27] $end
$var wire 1 TG c2 [26] $end
$var wire 1 UG c2 [25] $end
$var wire 1 VG c2 [24] $end
$var wire 1 WG c2 [23] $end
$var wire 1 XG c2 [22] $end
$var wire 1 YG c2 [21] $end
$var wire 1 ZG c2 [20] $end
$var wire 1 [G c2 [19] $end
$var wire 1 \G c2 [18] $end
$var wire 1 ]G c2 [17] $end
$var wire 1 ^G c2 [16] $end
$var wire 1 _G c2 [15] $end
$var wire 1 `G c2 [14] $end
$var wire 1 aG c2 [13] $end
$var wire 1 bG c2 [12] $end
$var wire 1 cG c2 [11] $end
$var wire 1 dG c2 [10] $end
$var wire 1 eG c2 [9] $end
$var wire 1 fG c2 [8] $end
$var wire 1 gG c2 [7] $end
$var wire 1 hG c2 [6] $end
$var wire 1 iG c2 [5] $end
$var wire 1 jG c2 [4] $end
$var wire 1 kG c2 [3] $end
$var wire 1 lG c2 [2] $end
$var wire 1 mG c2 [1] $end
$var wire 1 nG c2 [0] $end
$var wire 1 oG s [54] $end
$var wire 1 pG s [53] $end
$var wire 1 qG s [52] $end
$var wire 1 rG s [51] $end
$var wire 1 sG s [50] $end
$var wire 1 tG s [49] $end
$var wire 1 uG s [48] $end
$var wire 1 vG s [47] $end
$var wire 1 wG s [46] $end
$var wire 1 xG s [45] $end
$var wire 1 yG s [44] $end
$var wire 1 zG s [43] $end
$var wire 1 {G s [42] $end
$var wire 1 |G s [41] $end
$var wire 1 }G s [40] $end
$var wire 1 ~G s [39] $end
$var wire 1 !H s [38] $end
$var wire 1 "H s [37] $end
$var wire 1 #H s [36] $end
$var wire 1 $H s [35] $end
$var wire 1 %H s [34] $end
$var wire 1 &H s [33] $end
$var wire 1 'H s [32] $end
$var wire 1 (H s [31] $end
$var wire 1 )H s [30] $end
$var wire 1 *H s [29] $end
$var wire 1 +H s [28] $end
$var wire 1 ,H s [27] $end
$var wire 1 -H s [26] $end
$var wire 1 .H s [25] $end
$var wire 1 /H s [24] $end
$var wire 1 0H s [23] $end
$var wire 1 1H s [22] $end
$var wire 1 2H s [21] $end
$var wire 1 3H s [20] $end
$var wire 1 4H s [19] $end
$var wire 1 5H s [18] $end
$var wire 1 6H s [17] $end
$var wire 1 7H s [16] $end
$var wire 1 8H s [15] $end
$var wire 1 9H s [14] $end
$var wire 1 :H s [13] $end
$var wire 1 ;H s [12] $end
$var wire 1 <H s [11] $end
$var wire 1 =H s [10] $end
$var wire 1 >H s [9] $end
$var wire 1 ?H s [8] $end
$var wire 1 @H s [7] $end
$var wire 1 AH s [6] $end
$var wire 1 BH s [5] $end
$var wire 1 CH s [4] $end
$var wire 1 DH s [3] $end
$var wire 1 EH s [2] $end
$var wire 1 FH s [1] $end
$var wire 1 GH s [0] $end
$var wire 1 HH ca [54] $end
$var wire 1 IH ca [53] $end
$var wire 1 JH ca [52] $end
$var wire 1 KH ca [51] $end
$var wire 1 LH ca [50] $end
$var wire 1 MH ca [49] $end
$var wire 1 NH ca [48] $end
$var wire 1 OH ca [47] $end
$var wire 1 PH ca [46] $end
$var wire 1 QH ca [45] $end
$var wire 1 RH ca [44] $end
$var wire 1 SH ca [43] $end
$var wire 1 TH ca [42] $end
$var wire 1 UH ca [41] $end
$var wire 1 VH ca [40] $end
$var wire 1 WH ca [39] $end
$var wire 1 XH ca [38] $end
$var wire 1 YH ca [37] $end
$var wire 1 ZH ca [36] $end
$var wire 1 [H ca [35] $end
$var wire 1 \H ca [34] $end
$var wire 1 ]H ca [33] $end
$var wire 1 ^H ca [32] $end
$var wire 1 _H ca [31] $end
$var wire 1 `H ca [30] $end
$var wire 1 aH ca [29] $end
$var wire 1 bH ca [28] $end
$var wire 1 cH ca [27] $end
$var wire 1 dH ca [26] $end
$var wire 1 eH ca [25] $end
$var wire 1 fH ca [24] $end
$var wire 1 gH ca [23] $end
$var wire 1 hH ca [22] $end
$var wire 1 iH ca [21] $end
$var wire 1 jH ca [20] $end
$var wire 1 kH ca [19] $end
$var wire 1 lH ca [18] $end
$var wire 1 mH ca [17] $end
$var wire 1 nH ca [16] $end
$var wire 1 oH ca [15] $end
$var wire 1 pH ca [14] $end
$var wire 1 qH ca [13] $end
$var wire 1 rH ca [12] $end
$var wire 1 sH ca [11] $end
$var wire 1 tH ca [10] $end
$var wire 1 uH ca [9] $end
$var wire 1 vH ca [8] $end
$var wire 1 wH ca [7] $end
$var wire 1 xH ca [6] $end
$var wire 1 yH ca [5] $end
$var wire 1 zH ca [4] $end
$var wire 1 {H ca [3] $end
$var wire 1 |H ca [2] $end
$var wire 1 }H ca [1] $end
$var wire 1 ~H ca [0] $end
$upscope $end

$scope module l3_2 $end
$var parameter 32 AV size $end
$var wire 1 !I c0 [54] $end
$var wire 1 "I c0 [53] $end
$var wire 1 #I c0 [52] $end
$var wire 1 $I c0 [51] $end
$var wire 1 %I c0 [50] $end
$var wire 1 &I c0 [49] $end
$var wire 1 'I c0 [48] $end
$var wire 1 (I c0 [47] $end
$var wire 1 )I c0 [46] $end
$var wire 1 *I c0 [45] $end
$var wire 1 +I c0 [44] $end
$var wire 1 ,I c0 [43] $end
$var wire 1 -I c0 [42] $end
$var wire 1 .I c0 [41] $end
$var wire 1 /I c0 [40] $end
$var wire 1 0I c0 [39] $end
$var wire 1 1I c0 [38] $end
$var wire 1 2I c0 [37] $end
$var wire 1 3I c0 [36] $end
$var wire 1 4I c0 [35] $end
$var wire 1 5I c0 [34] $end
$var wire 1 6I c0 [33] $end
$var wire 1 7I c0 [32] $end
$var wire 1 8I c0 [31] $end
$var wire 1 9I c0 [30] $end
$var wire 1 :I c0 [29] $end
$var wire 1 ;I c0 [28] $end
$var wire 1 <I c0 [27] $end
$var wire 1 =I c0 [26] $end
$var wire 1 >I c0 [25] $end
$var wire 1 ?I c0 [24] $end
$var wire 1 @I c0 [23] $end
$var wire 1 AI c0 [22] $end
$var wire 1 BI c0 [21] $end
$var wire 1 CI c0 [20] $end
$var wire 1 DI c0 [19] $end
$var wire 1 EI c0 [18] $end
$var wire 1 FI c0 [17] $end
$var wire 1 GI c0 [16] $end
$var wire 1 HI c0 [15] $end
$var wire 1 II c0 [14] $end
$var wire 1 JI c0 [13] $end
$var wire 1 KI c0 [12] $end
$var wire 1 LI c0 [11] $end
$var wire 1 MI c0 [10] $end
$var wire 1 NI c0 [9] $end
$var wire 1 OI c0 [8] $end
$var wire 1 PI c0 [7] $end
$var wire 1 QI c0 [6] $end
$var wire 1 RI c0 [5] $end
$var wire 1 SI c0 [4] $end
$var wire 1 TI c0 [3] $end
$var wire 1 UI c0 [2] $end
$var wire 1 VI c0 [1] $end
$var wire 1 WI c0 [0] $end
$var wire 1 XI c1 [54] $end
$var wire 1 YI c1 [53] $end
$var wire 1 ZI c1 [52] $end
$var wire 1 [I c1 [51] $end
$var wire 1 \I c1 [50] $end
$var wire 1 ]I c1 [49] $end
$var wire 1 ^I c1 [48] $end
$var wire 1 _I c1 [47] $end
$var wire 1 `I c1 [46] $end
$var wire 1 aI c1 [45] $end
$var wire 1 bI c1 [44] $end
$var wire 1 cI c1 [43] $end
$var wire 1 dI c1 [42] $end
$var wire 1 eI c1 [41] $end
$var wire 1 fI c1 [40] $end
$var wire 1 gI c1 [39] $end
$var wire 1 hI c1 [38] $end
$var wire 1 iI c1 [37] $end
$var wire 1 jI c1 [36] $end
$var wire 1 kI c1 [35] $end
$var wire 1 lI c1 [34] $end
$var wire 1 mI c1 [33] $end
$var wire 1 nI c1 [32] $end
$var wire 1 oI c1 [31] $end
$var wire 1 pI c1 [30] $end
$var wire 1 qI c1 [29] $end
$var wire 1 rI c1 [28] $end
$var wire 1 sI c1 [27] $end
$var wire 1 tI c1 [26] $end
$var wire 1 uI c1 [25] $end
$var wire 1 vI c1 [24] $end
$var wire 1 wI c1 [23] $end
$var wire 1 xI c1 [22] $end
$var wire 1 yI c1 [21] $end
$var wire 1 zI c1 [20] $end
$var wire 1 {I c1 [19] $end
$var wire 1 |I c1 [18] $end
$var wire 1 }I c1 [17] $end
$var wire 1 ~I c1 [16] $end
$var wire 1 !J c1 [15] $end
$var wire 1 "J c1 [14] $end
$var wire 1 #J c1 [13] $end
$var wire 1 $J c1 [12] $end
$var wire 1 %J c1 [11] $end
$var wire 1 &J c1 [10] $end
$var wire 1 'J c1 [9] $end
$var wire 1 (J c1 [8] $end
$var wire 1 )J c1 [7] $end
$var wire 1 *J c1 [6] $end
$var wire 1 +J c1 [5] $end
$var wire 1 ,J c1 [4] $end
$var wire 1 -J c1 [3] $end
$var wire 1 .J c1 [2] $end
$var wire 1 /J c1 [1] $end
$var wire 1 0J c1 [0] $end
$var wire 1 1J c2 [54] $end
$var wire 1 2J c2 [53] $end
$var wire 1 3J c2 [52] $end
$var wire 1 4J c2 [51] $end
$var wire 1 5J c2 [50] $end
$var wire 1 6J c2 [49] $end
$var wire 1 7J c2 [48] $end
$var wire 1 8J c2 [47] $end
$var wire 1 9J c2 [46] $end
$var wire 1 :J c2 [45] $end
$var wire 1 ;J c2 [44] $end
$var wire 1 <J c2 [43] $end
$var wire 1 =J c2 [42] $end
$var wire 1 >J c2 [41] $end
$var wire 1 ?J c2 [40] $end
$var wire 1 @J c2 [39] $end
$var wire 1 AJ c2 [38] $end
$var wire 1 BJ c2 [37] $end
$var wire 1 CJ c2 [36] $end
$var wire 1 DJ c2 [35] $end
$var wire 1 EJ c2 [34] $end
$var wire 1 FJ c2 [33] $end
$var wire 1 GJ c2 [32] $end
$var wire 1 HJ c2 [31] $end
$var wire 1 IJ c2 [30] $end
$var wire 1 JJ c2 [29] $end
$var wire 1 KJ c2 [28] $end
$var wire 1 LJ c2 [27] $end
$var wire 1 MJ c2 [26] $end
$var wire 1 NJ c2 [25] $end
$var wire 1 OJ c2 [24] $end
$var wire 1 PJ c2 [23] $end
$var wire 1 QJ c2 [22] $end
$var wire 1 RJ c2 [21] $end
$var wire 1 SJ c2 [20] $end
$var wire 1 TJ c2 [19] $end
$var wire 1 UJ c2 [18] $end
$var wire 1 VJ c2 [17] $end
$var wire 1 WJ c2 [16] $end
$var wire 1 XJ c2 [15] $end
$var wire 1 YJ c2 [14] $end
$var wire 1 ZJ c2 [13] $end
$var wire 1 [J c2 [12] $end
$var wire 1 \J c2 [11] $end
$var wire 1 ]J c2 [10] $end
$var wire 1 ^J c2 [9] $end
$var wire 1 _J c2 [8] $end
$var wire 1 `J c2 [7] $end
$var wire 1 aJ c2 [6] $end
$var wire 1 bJ c2 [5] $end
$var wire 1 cJ c2 [4] $end
$var wire 1 dJ c2 [3] $end
$var wire 1 eJ c2 [2] $end
$var wire 1 fJ c2 [1] $end
$var wire 1 gJ c2 [0] $end
$var wire 1 hJ s [54] $end
$var wire 1 iJ s [53] $end
$var wire 1 jJ s [52] $end
$var wire 1 kJ s [51] $end
$var wire 1 lJ s [50] $end
$var wire 1 mJ s [49] $end
$var wire 1 nJ s [48] $end
$var wire 1 oJ s [47] $end
$var wire 1 pJ s [46] $end
$var wire 1 qJ s [45] $end
$var wire 1 rJ s [44] $end
$var wire 1 sJ s [43] $end
$var wire 1 tJ s [42] $end
$var wire 1 uJ s [41] $end
$var wire 1 vJ s [40] $end
$var wire 1 wJ s [39] $end
$var wire 1 xJ s [38] $end
$var wire 1 yJ s [37] $end
$var wire 1 zJ s [36] $end
$var wire 1 {J s [35] $end
$var wire 1 |J s [34] $end
$var wire 1 }J s [33] $end
$var wire 1 ~J s [32] $end
$var wire 1 !K s [31] $end
$var wire 1 "K s [30] $end
$var wire 1 #K s [29] $end
$var wire 1 $K s [28] $end
$var wire 1 %K s [27] $end
$var wire 1 &K s [26] $end
$var wire 1 'K s [25] $end
$var wire 1 (K s [24] $end
$var wire 1 )K s [23] $end
$var wire 1 *K s [22] $end
$var wire 1 +K s [21] $end
$var wire 1 ,K s [20] $end
$var wire 1 -K s [19] $end
$var wire 1 .K s [18] $end
$var wire 1 /K s [17] $end
$var wire 1 0K s [16] $end
$var wire 1 1K s [15] $end
$var wire 1 2K s [14] $end
$var wire 1 3K s [13] $end
$var wire 1 4K s [12] $end
$var wire 1 5K s [11] $end
$var wire 1 6K s [10] $end
$var wire 1 7K s [9] $end
$var wire 1 8K s [8] $end
$var wire 1 9K s [7] $end
$var wire 1 :K s [6] $end
$var wire 1 ;K s [5] $end
$var wire 1 <K s [4] $end
$var wire 1 =K s [3] $end
$var wire 1 >K s [2] $end
$var wire 1 ?K s [1] $end
$var wire 1 @K s [0] $end
$var wire 1 AK ca [54] $end
$var wire 1 BK ca [53] $end
$var wire 1 CK ca [52] $end
$var wire 1 DK ca [51] $end
$var wire 1 EK ca [50] $end
$var wire 1 FK ca [49] $end
$var wire 1 GK ca [48] $end
$var wire 1 HK ca [47] $end
$var wire 1 IK ca [46] $end
$var wire 1 JK ca [45] $end
$var wire 1 KK ca [44] $end
$var wire 1 LK ca [43] $end
$var wire 1 MK ca [42] $end
$var wire 1 NK ca [41] $end
$var wire 1 OK ca [40] $end
$var wire 1 PK ca [39] $end
$var wire 1 QK ca [38] $end
$var wire 1 RK ca [37] $end
$var wire 1 SK ca [36] $end
$var wire 1 TK ca [35] $end
$var wire 1 UK ca [34] $end
$var wire 1 VK ca [33] $end
$var wire 1 WK ca [32] $end
$var wire 1 XK ca [31] $end
$var wire 1 YK ca [30] $end
$var wire 1 ZK ca [29] $end
$var wire 1 [K ca [28] $end
$var wire 1 \K ca [27] $end
$var wire 1 ]K ca [26] $end
$var wire 1 ^K ca [25] $end
$var wire 1 _K ca [24] $end
$var wire 1 `K ca [23] $end
$var wire 1 aK ca [22] $end
$var wire 1 bK ca [21] $end
$var wire 1 cK ca [20] $end
$var wire 1 dK ca [19] $end
$var wire 1 eK ca [18] $end
$var wire 1 fK ca [17] $end
$var wire 1 gK ca [16] $end
$var wire 1 hK ca [15] $end
$var wire 1 iK ca [14] $end
$var wire 1 jK ca [13] $end
$var wire 1 kK ca [12] $end
$var wire 1 lK ca [11] $end
$var wire 1 mK ca [10] $end
$var wire 1 nK ca [9] $end
$var wire 1 oK ca [8] $end
$var wire 1 pK ca [7] $end
$var wire 1 qK ca [6] $end
$var wire 1 rK ca [5] $end
$var wire 1 sK ca [4] $end
$var wire 1 tK ca [3] $end
$var wire 1 uK ca [2] $end
$var wire 1 vK ca [1] $end
$var wire 1 wK ca [0] $end
$upscope $end

$scope module l4 $end
$var parameter 32 BV size $end
$var wire 1 CV p1 [63] $end
$var wire 1 DV p1 [62] $end
$var wire 1 EV p1 [61] $end
$var wire 1 FV p1 [60] $end
$var wire 1 GV p1 [59] $end
$var wire 1 HV p1 [58] $end
$var wire 1 IV p1 [57] $end
$var wire 1 JV p1 [56] $end
$var wire 1 KV p1 [55] $end
$var wire 1 LV p1 [54] $end
$var wire 1 MV p1 [53] $end
$var wire 1 NV p1 [52] $end
$var wire 1 OV p1 [51] $end
$var wire 1 PV p1 [50] $end
$var wire 1 QV p1 [49] $end
$var wire 1 RV p1 [48] $end
$var wire 1 SV p1 [47] $end
$var wire 1 TV p1 [46] $end
$var wire 1 UV p1 [45] $end
$var wire 1 VV p1 [44] $end
$var wire 1 WV p1 [43] $end
$var wire 1 XV p1 [42] $end
$var wire 1 YV p1 [41] $end
$var wire 1 ZV p1 [40] $end
$var wire 1 [V p1 [39] $end
$var wire 1 \V p1 [38] $end
$var wire 1 ]V p1 [37] $end
$var wire 1 ^V p1 [36] $end
$var wire 1 _V p1 [35] $end
$var wire 1 `V p1 [34] $end
$var wire 1 aV p1 [33] $end
$var wire 1 bV p1 [32] $end
$var wire 1 cV p1 [31] $end
$var wire 1 dV p1 [30] $end
$var wire 1 eV p1 [29] $end
$var wire 1 fV p1 [28] $end
$var wire 1 gV p1 [27] $end
$var wire 1 hV p1 [26] $end
$var wire 1 iV p1 [25] $end
$var wire 1 jV p1 [24] $end
$var wire 1 kV p1 [23] $end
$var wire 1 lV p1 [22] $end
$var wire 1 mV p1 [21] $end
$var wire 1 nV p1 [20] $end
$var wire 1 oV p1 [19] $end
$var wire 1 pV p1 [18] $end
$var wire 1 qV p1 [17] $end
$var wire 1 rV p1 [16] $end
$var wire 1 sV p1 [15] $end
$var wire 1 tV p1 [14] $end
$var wire 1 uV p1 [13] $end
$var wire 1 vV p1 [12] $end
$var wire 1 wV p1 [11] $end
$var wire 1 xV p1 [10] $end
$var wire 1 yV p1 [9] $end
$var wire 1 zV p1 [8] $end
$var wire 1 {V p1 [7] $end
$var wire 1 |V p1 [6] $end
$var wire 1 }V p1 [5] $end
$var wire 1 ~V p1 [4] $end
$var wire 1 !W p1 [3] $end
$var wire 1 "W p1 [2] $end
$var wire 1 #W p1 [1] $end
$var wire 1 $W p1 [0] $end
$var wire 1 %W p2 [63] $end
$var wire 1 &W p2 [62] $end
$var wire 1 'W p2 [61] $end
$var wire 1 (W p2 [60] $end
$var wire 1 )W p2 [59] $end
$var wire 1 *W p2 [58] $end
$var wire 1 +W p2 [57] $end
$var wire 1 ,W p2 [56] $end
$var wire 1 -W p2 [55] $end
$var wire 1 .W p2 [54] $end
$var wire 1 /W p2 [53] $end
$var wire 1 0W p2 [52] $end
$var wire 1 1W p2 [51] $end
$var wire 1 2W p2 [50] $end
$var wire 1 3W p2 [49] $end
$var wire 1 4W p2 [48] $end
$var wire 1 5W p2 [47] $end
$var wire 1 6W p2 [46] $end
$var wire 1 7W p2 [45] $end
$var wire 1 8W p2 [44] $end
$var wire 1 9W p2 [43] $end
$var wire 1 :W p2 [42] $end
$var wire 1 ;W p2 [41] $end
$var wire 1 <W p2 [40] $end
$var wire 1 =W p2 [39] $end
$var wire 1 >W p2 [38] $end
$var wire 1 ?W p2 [37] $end
$var wire 1 @W p2 [36] $end
$var wire 1 AW p2 [35] $end
$var wire 1 BW p2 [34] $end
$var wire 1 CW p2 [33] $end
$var wire 1 DW p2 [32] $end
$var wire 1 EW p2 [31] $end
$var wire 1 FW p2 [30] $end
$var wire 1 GW p2 [29] $end
$var wire 1 HW p2 [28] $end
$var wire 1 IW p2 [27] $end
$var wire 1 JW p2 [26] $end
$var wire 1 KW p2 [25] $end
$var wire 1 LW p2 [24] $end
$var wire 1 MW p2 [23] $end
$var wire 1 NW p2 [22] $end
$var wire 1 OW p2 [21] $end
$var wire 1 PW p2 [20] $end
$var wire 1 QW p2 [19] $end
$var wire 1 RW p2 [18] $end
$var wire 1 SW p2 [17] $end
$var wire 1 TW p2 [16] $end
$var wire 1 UW p2 [15] $end
$var wire 1 VW p2 [14] $end
$var wire 1 WW p2 [13] $end
$var wire 1 XW p2 [12] $end
$var wire 1 YW p2 [11] $end
$var wire 1 ZW p2 [10] $end
$var wire 1 [W p2 [9] $end
$var wire 1 \W p2 [8] $end
$var wire 1 ]W p2 [7] $end
$var wire 1 ^W p2 [6] $end
$var wire 1 _W p2 [5] $end
$var wire 1 `W p2 [4] $end
$var wire 1 aW p2 [3] $end
$var wire 1 bW p2 [2] $end
$var wire 1 cW p2 [1] $end
$var wire 1 dW p2 [0] $end
$var wire 1 eW p3 [63] $end
$var wire 1 fW p3 [62] $end
$var wire 1 gW p3 [61] $end
$var wire 1 hW p3 [60] $end
$var wire 1 iW p3 [59] $end
$var wire 1 jW p3 [58] $end
$var wire 1 kW p3 [57] $end
$var wire 1 lW p3 [56] $end
$var wire 1 mW p3 [55] $end
$var wire 1 nW p3 [54] $end
$var wire 1 oW p3 [53] $end
$var wire 1 pW p3 [52] $end
$var wire 1 qW p3 [51] $end
$var wire 1 rW p3 [50] $end
$var wire 1 sW p3 [49] $end
$var wire 1 tW p3 [48] $end
$var wire 1 uW p3 [47] $end
$var wire 1 vW p3 [46] $end
$var wire 1 wW p3 [45] $end
$var wire 1 xW p3 [44] $end
$var wire 1 yW p3 [43] $end
$var wire 1 zW p3 [42] $end
$var wire 1 {W p3 [41] $end
$var wire 1 |W p3 [40] $end
$var wire 1 }W p3 [39] $end
$var wire 1 ~W p3 [38] $end
$var wire 1 !X p3 [37] $end
$var wire 1 "X p3 [36] $end
$var wire 1 #X p3 [35] $end
$var wire 1 $X p3 [34] $end
$var wire 1 %X p3 [33] $end
$var wire 1 &X p3 [32] $end
$var wire 1 'X p3 [31] $end
$var wire 1 (X p3 [30] $end
$var wire 1 )X p3 [29] $end
$var wire 1 *X p3 [28] $end
$var wire 1 +X p3 [27] $end
$var wire 1 ,X p3 [26] $end
$var wire 1 -X p3 [25] $end
$var wire 1 .X p3 [24] $end
$var wire 1 /X p3 [23] $end
$var wire 1 0X p3 [22] $end
$var wire 1 1X p3 [21] $end
$var wire 1 2X p3 [20] $end
$var wire 1 3X p3 [19] $end
$var wire 1 4X p3 [18] $end
$var wire 1 5X p3 [17] $end
$var wire 1 6X p3 [16] $end
$var wire 1 7X p3 [15] $end
$var wire 1 8X p3 [14] $end
$var wire 1 9X p3 [13] $end
$var wire 1 :X p3 [12] $end
$var wire 1 ;X p3 [11] $end
$var wire 1 <X p3 [10] $end
$var wire 1 =X p3 [9] $end
$var wire 1 >X p3 [8] $end
$var wire 1 ?X p3 [7] $end
$var wire 1 @X p3 [6] $end
$var wire 1 AX p3 [5] $end
$var wire 1 BX p3 [4] $end
$var wire 1 CX p3 [3] $end
$var wire 1 DX p3 [2] $end
$var wire 1 EX p3 [1] $end
$var wire 1 FX p3 [0] $end
$var wire 1 |K c1 [63] $end
$var wire 1 }K c1 [62] $end
$var wire 1 ~K c1 [61] $end
$var wire 1 !L c1 [60] $end
$var wire 1 "L c1 [59] $end
$var wire 1 #L c1 [58] $end
$var wire 1 $L c1 [57] $end
$var wire 1 %L c1 [56] $end
$var wire 1 &L c1 [55] $end
$var wire 1 'L c1 [54] $end
$var wire 1 (L c1 [53] $end
$var wire 1 )L c1 [52] $end
$var wire 1 *L c1 [51] $end
$var wire 1 +L c1 [50] $end
$var wire 1 ,L c1 [49] $end
$var wire 1 -L c1 [48] $end
$var wire 1 .L c1 [47] $end
$var wire 1 /L c1 [46] $end
$var wire 1 0L c1 [45] $end
$var wire 1 1L c1 [44] $end
$var wire 1 2L c1 [43] $end
$var wire 1 3L c1 [42] $end
$var wire 1 4L c1 [41] $end
$var wire 1 5L c1 [40] $end
$var wire 1 6L c1 [39] $end
$var wire 1 7L c1 [38] $end
$var wire 1 8L c1 [37] $end
$var wire 1 9L c1 [36] $end
$var wire 1 :L c1 [35] $end
$var wire 1 ;L c1 [34] $end
$var wire 1 <L c1 [33] $end
$var wire 1 =L c1 [32] $end
$var wire 1 >L c1 [31] $end
$var wire 1 ?L c1 [30] $end
$var wire 1 @L c1 [29] $end
$var wire 1 AL c1 [28] $end
$var wire 1 BL c1 [27] $end
$var wire 1 CL c1 [26] $end
$var wire 1 DL c1 [25] $end
$var wire 1 EL c1 [24] $end
$var wire 1 FL c1 [23] $end
$var wire 1 GL c1 [22] $end
$var wire 1 HL c1 [21] $end
$var wire 1 IL c1 [20] $end
$var wire 1 JL c1 [19] $end
$var wire 1 KL c1 [18] $end
$var wire 1 LL c1 [17] $end
$var wire 1 ML c1 [16] $end
$var wire 1 NL c1 [15] $end
$var wire 1 OL c1 [14] $end
$var wire 1 PL c1 [13] $end
$var wire 1 QL c1 [12] $end
$var wire 1 RL c1 [11] $end
$var wire 1 SL c1 [10] $end
$var wire 1 TL c1 [9] $end
$var wire 1 UL c1 [8] $end
$var wire 1 VL c1 [7] $end
$var wire 1 WL c1 [6] $end
$var wire 1 XL c1 [5] $end
$var wire 1 YL c1 [4] $end
$var wire 1 ZL c1 [3] $end
$var wire 1 [L c1 [2] $end
$var wire 1 \L c1 [1] $end
$var wire 1 ]L c1 [0] $end
$var wire 1 ^L c2 [63] $end
$var wire 1 _L c2 [62] $end
$var wire 1 `L c2 [61] $end
$var wire 1 aL c2 [60] $end
$var wire 1 bL c2 [59] $end
$var wire 1 cL c2 [58] $end
$var wire 1 dL c2 [57] $end
$var wire 1 eL c2 [56] $end
$var wire 1 fL c2 [55] $end
$var wire 1 gL c2 [54] $end
$var wire 1 hL c2 [53] $end
$var wire 1 iL c2 [52] $end
$var wire 1 jL c2 [51] $end
$var wire 1 kL c2 [50] $end
$var wire 1 lL c2 [49] $end
$var wire 1 mL c2 [48] $end
$var wire 1 nL c2 [47] $end
$var wire 1 oL c2 [46] $end
$var wire 1 pL c2 [45] $end
$var wire 1 qL c2 [44] $end
$var wire 1 rL c2 [43] $end
$var wire 1 sL c2 [42] $end
$var wire 1 tL c2 [41] $end
$var wire 1 uL c2 [40] $end
$var wire 1 vL c2 [39] $end
$var wire 1 wL c2 [38] $end
$var wire 1 xL c2 [37] $end
$var wire 1 yL c2 [36] $end
$var wire 1 zL c2 [35] $end
$var wire 1 {L c2 [34] $end
$var wire 1 |L c2 [33] $end
$var wire 1 }L c2 [32] $end
$var wire 1 ~L c2 [31] $end
$var wire 1 !M c2 [30] $end
$var wire 1 "M c2 [29] $end
$var wire 1 #M c2 [28] $end
$var wire 1 $M c2 [27] $end
$var wire 1 %M c2 [26] $end
$var wire 1 &M c2 [25] $end
$var wire 1 'M c2 [24] $end
$var wire 1 (M c2 [23] $end
$var wire 1 )M c2 [22] $end
$var wire 1 *M c2 [21] $end
$var wire 1 +M c2 [20] $end
$var wire 1 ,M c2 [19] $end
$var wire 1 -M c2 [18] $end
$var wire 1 .M c2 [17] $end
$var wire 1 /M c2 [16] $end
$var wire 1 0M c2 [15] $end
$var wire 1 1M c2 [14] $end
$var wire 1 2M c2 [13] $end
$var wire 1 3M c2 [12] $end
$var wire 1 4M c2 [11] $end
$var wire 1 5M c2 [10] $end
$var wire 1 6M c2 [9] $end
$var wire 1 7M c2 [8] $end
$var wire 1 8M c2 [7] $end
$var wire 1 9M c2 [6] $end
$var wire 1 :M c2 [5] $end
$var wire 1 ;M c2 [4] $end
$var wire 1 <M c2 [3] $end
$var wire 1 =M c2 [2] $end
$var wire 1 >M c2 [1] $end
$var wire 1 ?M c2 [0] $end
$var wire 1 @M c3 [63] $end
$var wire 1 AM c3 [62] $end
$var wire 1 BM c3 [61] $end
$var wire 1 CM c3 [60] $end
$var wire 1 DM c3 [59] $end
$var wire 1 EM c3 [58] $end
$var wire 1 FM c3 [57] $end
$var wire 1 GM c3 [56] $end
$var wire 1 HM c3 [55] $end
$var wire 1 IM c3 [54] $end
$var wire 1 JM c3 [53] $end
$var wire 1 KM c3 [52] $end
$var wire 1 LM c3 [51] $end
$var wire 1 MM c3 [50] $end
$var wire 1 NM c3 [49] $end
$var wire 1 OM c3 [48] $end
$var wire 1 PM c3 [47] $end
$var wire 1 QM c3 [46] $end
$var wire 1 RM c3 [45] $end
$var wire 1 SM c3 [44] $end
$var wire 1 TM c3 [43] $end
$var wire 1 UM c3 [42] $end
$var wire 1 VM c3 [41] $end
$var wire 1 WM c3 [40] $end
$var wire 1 XM c3 [39] $end
$var wire 1 YM c3 [38] $end
$var wire 1 ZM c3 [37] $end
$var wire 1 [M c3 [36] $end
$var wire 1 \M c3 [35] $end
$var wire 1 ]M c3 [34] $end
$var wire 1 ^M c3 [33] $end
$var wire 1 _M c3 [32] $end
$var wire 1 `M c3 [31] $end
$var wire 1 aM c3 [30] $end
$var wire 1 bM c3 [29] $end
$var wire 1 cM c3 [28] $end
$var wire 1 dM c3 [27] $end
$var wire 1 eM c3 [26] $end
$var wire 1 fM c3 [25] $end
$var wire 1 gM c3 [24] $end
$var wire 1 hM c3 [23] $end
$var wire 1 iM c3 [22] $end
$var wire 1 jM c3 [21] $end
$var wire 1 kM c3 [20] $end
$var wire 1 lM c3 [19] $end
$var wire 1 mM c3 [18] $end
$var wire 1 nM c3 [17] $end
$var wire 1 oM c3 [16] $end
$var wire 1 pM c3 [15] $end
$var wire 1 qM c3 [14] $end
$var wire 1 rM c3 [13] $end
$var wire 1 sM c3 [12] $end
$var wire 1 tM c3 [11] $end
$var wire 1 uM c3 [10] $end
$var wire 1 vM c3 [9] $end
$var wire 1 wM c3 [8] $end
$var wire 1 xM c3 [7] $end
$var wire 1 yM c3 [6] $end
$var wire 1 zM c3 [5] $end
$var wire 1 {M c3 [4] $end
$var wire 1 |M c3 [3] $end
$var wire 1 }M c3 [2] $end
$var wire 1 ~M c3 [1] $end
$var wire 1 !N c3 [0] $end
$var wire 1 "N c4 [63] $end
$var wire 1 #N c4 [62] $end
$var wire 1 $N c4 [61] $end
$var wire 1 %N c4 [60] $end
$var wire 1 &N c4 [59] $end
$var wire 1 'N c4 [58] $end
$var wire 1 (N c4 [57] $end
$var wire 1 )N c4 [56] $end
$var wire 1 *N c4 [55] $end
$var wire 1 +N c4 [54] $end
$var wire 1 ,N c4 [53] $end
$var wire 1 -N c4 [52] $end
$var wire 1 .N c4 [51] $end
$var wire 1 /N c4 [50] $end
$var wire 1 0N c4 [49] $end
$var wire 1 1N c4 [48] $end
$var wire 1 2N c4 [47] $end
$var wire 1 3N c4 [46] $end
$var wire 1 4N c4 [45] $end
$var wire 1 5N c4 [44] $end
$var wire 1 6N c4 [43] $end
$var wire 1 7N c4 [42] $end
$var wire 1 8N c4 [41] $end
$var wire 1 9N c4 [40] $end
$var wire 1 :N c4 [39] $end
$var wire 1 ;N c4 [38] $end
$var wire 1 <N c4 [37] $end
$var wire 1 =N c4 [36] $end
$var wire 1 >N c4 [35] $end
$var wire 1 ?N c4 [34] $end
$var wire 1 @N c4 [33] $end
$var wire 1 AN c4 [32] $end
$var wire 1 BN c4 [31] $end
$var wire 1 CN c4 [30] $end
$var wire 1 DN c4 [29] $end
$var wire 1 EN c4 [28] $end
$var wire 1 FN c4 [27] $end
$var wire 1 GN c4 [26] $end
$var wire 1 HN c4 [25] $end
$var wire 1 IN c4 [24] $end
$var wire 1 JN c4 [23] $end
$var wire 1 KN c4 [22] $end
$var wire 1 LN c4 [21] $end
$var wire 1 MN c4 [20] $end
$var wire 1 NN c4 [19] $end
$var wire 1 ON c4 [18] $end
$var wire 1 PN c4 [17] $end
$var wire 1 QN c4 [16] $end
$var wire 1 RN c4 [15] $end
$var wire 1 SN c4 [14] $end
$var wire 1 TN c4 [13] $end
$var wire 1 UN c4 [12] $end
$var wire 1 VN c4 [11] $end
$var wire 1 WN c4 [10] $end
$var wire 1 XN c4 [9] $end
$var wire 1 YN c4 [8] $end
$var wire 1 ZN c4 [7] $end
$var wire 1 [N c4 [6] $end
$var wire 1 \N c4 [5] $end
$var wire 1 ]N c4 [4] $end
$var wire 1 ^N c4 [3] $end
$var wire 1 _N c4 [2] $end
$var wire 1 `N c4 [1] $end
$var wire 1 aN c4 [0] $end
$var wire 1 &P cin [63] $end
$var wire 1 'P cin [62] $end
$var wire 1 (P cin [61] $end
$var wire 1 )P cin [60] $end
$var wire 1 *P cin [59] $end
$var wire 1 +P cin [58] $end
$var wire 1 ,P cin [57] $end
$var wire 1 -P cin [56] $end
$var wire 1 .P cin [55] $end
$var wire 1 /P cin [54] $end
$var wire 1 0P cin [53] $end
$var wire 1 1P cin [52] $end
$var wire 1 2P cin [51] $end
$var wire 1 3P cin [50] $end
$var wire 1 4P cin [49] $end
$var wire 1 5P cin [48] $end
$var wire 1 6P cin [47] $end
$var wire 1 7P cin [46] $end
$var wire 1 8P cin [45] $end
$var wire 1 9P cin [44] $end
$var wire 1 :P cin [43] $end
$var wire 1 ;P cin [42] $end
$var wire 1 <P cin [41] $end
$var wire 1 =P cin [40] $end
$var wire 1 >P cin [39] $end
$var wire 1 ?P cin [38] $end
$var wire 1 @P cin [37] $end
$var wire 1 AP cin [36] $end
$var wire 1 BP cin [35] $end
$var wire 1 CP cin [34] $end
$var wire 1 DP cin [33] $end
$var wire 1 EP cin [32] $end
$var wire 1 FP cin [31] $end
$var wire 1 GP cin [30] $end
$var wire 1 HP cin [29] $end
$var wire 1 IP cin [28] $end
$var wire 1 JP cin [27] $end
$var wire 1 KP cin [26] $end
$var wire 1 LP cin [25] $end
$var wire 1 MP cin [24] $end
$var wire 1 NP cin [23] $end
$var wire 1 OP cin [22] $end
$var wire 1 PP cin [21] $end
$var wire 1 QP cin [20] $end
$var wire 1 RP cin [19] $end
$var wire 1 SP cin [18] $end
$var wire 1 TP cin [17] $end
$var wire 1 UP cin [16] $end
$var wire 1 VP cin [15] $end
$var wire 1 WP cin [14] $end
$var wire 1 XP cin [13] $end
$var wire 1 YP cin [12] $end
$var wire 1 ZP cin [11] $end
$var wire 1 [P cin [10] $end
$var wire 1 \P cin [9] $end
$var wire 1 ]P cin [8] $end
$var wire 1 ^P cin [7] $end
$var wire 1 _P cin [6] $end
$var wire 1 `P cin [5] $end
$var wire 1 aP cin [4] $end
$var wire 1 bP cin [3] $end
$var wire 1 cP cin [2] $end
$var wire 1 dP cin [1] $end
$var wire 1 eP cin [0] $end
$var wire 1 fP cout [63] $end
$var wire 1 gP cout [62] $end
$var wire 1 hP cout [61] $end
$var wire 1 iP cout [60] $end
$var wire 1 jP cout [59] $end
$var wire 1 kP cout [58] $end
$var wire 1 lP cout [57] $end
$var wire 1 mP cout [56] $end
$var wire 1 nP cout [55] $end
$var wire 1 oP cout [54] $end
$var wire 1 pP cout [53] $end
$var wire 1 qP cout [52] $end
$var wire 1 rP cout [51] $end
$var wire 1 sP cout [50] $end
$var wire 1 tP cout [49] $end
$var wire 1 uP cout [48] $end
$var wire 1 vP cout [47] $end
$var wire 1 wP cout [46] $end
$var wire 1 xP cout [45] $end
$var wire 1 yP cout [44] $end
$var wire 1 zP cout [43] $end
$var wire 1 {P cout [42] $end
$var wire 1 |P cout [41] $end
$var wire 1 }P cout [40] $end
$var wire 1 ~P cout [39] $end
$var wire 1 !Q cout [38] $end
$var wire 1 "Q cout [37] $end
$var wire 1 #Q cout [36] $end
$var wire 1 $Q cout [35] $end
$var wire 1 %Q cout [34] $end
$var wire 1 &Q cout [33] $end
$var wire 1 'Q cout [32] $end
$var wire 1 (Q cout [31] $end
$var wire 1 )Q cout [30] $end
$var wire 1 *Q cout [29] $end
$var wire 1 +Q cout [28] $end
$var wire 1 ,Q cout [27] $end
$var wire 1 -Q cout [26] $end
$var wire 1 .Q cout [25] $end
$var wire 1 /Q cout [24] $end
$var wire 1 0Q cout [23] $end
$var wire 1 1Q cout [22] $end
$var wire 1 2Q cout [21] $end
$var wire 1 3Q cout [20] $end
$var wire 1 4Q cout [19] $end
$var wire 1 5Q cout [18] $end
$var wire 1 6Q cout [17] $end
$var wire 1 7Q cout [16] $end
$var wire 1 8Q cout [15] $end
$var wire 1 9Q cout [14] $end
$var wire 1 :Q cout [13] $end
$var wire 1 ;Q cout [12] $end
$var wire 1 <Q cout [11] $end
$var wire 1 =Q cout [10] $end
$var wire 1 >Q cout [9] $end
$var wire 1 ?Q cout [8] $end
$var wire 1 @Q cout [7] $end
$var wire 1 AQ cout [6] $end
$var wire 1 BQ cout [5] $end
$var wire 1 CQ cout [4] $end
$var wire 1 DQ cout [3] $end
$var wire 1 EQ cout [2] $end
$var wire 1 FQ cout [1] $end
$var wire 1 GQ cout [0] $end
$var wire 1 bN s [63] $end
$var wire 1 cN s [62] $end
$var wire 1 dN s [61] $end
$var wire 1 eN s [60] $end
$var wire 1 fN s [59] $end
$var wire 1 gN s [58] $end
$var wire 1 hN s [57] $end
$var wire 1 iN s [56] $end
$var wire 1 jN s [55] $end
$var wire 1 kN s [54] $end
$var wire 1 lN s [53] $end
$var wire 1 mN s [52] $end
$var wire 1 nN s [51] $end
$var wire 1 oN s [50] $end
$var wire 1 pN s [49] $end
$var wire 1 qN s [48] $end
$var wire 1 rN s [47] $end
$var wire 1 sN s [46] $end
$var wire 1 tN s [45] $end
$var wire 1 uN s [44] $end
$var wire 1 vN s [43] $end
$var wire 1 wN s [42] $end
$var wire 1 xN s [41] $end
$var wire 1 yN s [40] $end
$var wire 1 zN s [39] $end
$var wire 1 {N s [38] $end
$var wire 1 |N s [37] $end
$var wire 1 }N s [36] $end
$var wire 1 ~N s [35] $end
$var wire 1 !O s [34] $end
$var wire 1 "O s [33] $end
$var wire 1 #O s [32] $end
$var wire 1 $O s [31] $end
$var wire 1 %O s [30] $end
$var wire 1 &O s [29] $end
$var wire 1 'O s [28] $end
$var wire 1 (O s [27] $end
$var wire 1 )O s [26] $end
$var wire 1 *O s [25] $end
$var wire 1 +O s [24] $end
$var wire 1 ,O s [23] $end
$var wire 1 -O s [22] $end
$var wire 1 .O s [21] $end
$var wire 1 /O s [20] $end
$var wire 1 0O s [19] $end
$var wire 1 1O s [18] $end
$var wire 1 2O s [17] $end
$var wire 1 3O s [16] $end
$var wire 1 4O s [15] $end
$var wire 1 5O s [14] $end
$var wire 1 6O s [13] $end
$var wire 1 7O s [12] $end
$var wire 1 8O s [11] $end
$var wire 1 9O s [10] $end
$var wire 1 :O s [9] $end
$var wire 1 ;O s [8] $end
$var wire 1 <O s [7] $end
$var wire 1 =O s [6] $end
$var wire 1 >O s [5] $end
$var wire 1 ?O s [4] $end
$var wire 1 @O s [3] $end
$var wire 1 AO s [2] $end
$var wire 1 BO s [1] $end
$var wire 1 CO s [0] $end
$var wire 1 DO ca [63] $end
$var wire 1 EO ca [62] $end
$var wire 1 FO ca [61] $end
$var wire 1 GO ca [60] $end
$var wire 1 HO ca [59] $end
$var wire 1 IO ca [58] $end
$var wire 1 JO ca [57] $end
$var wire 1 KO ca [56] $end
$var wire 1 LO ca [55] $end
$var wire 1 MO ca [54] $end
$var wire 1 NO ca [53] $end
$var wire 1 OO ca [52] $end
$var wire 1 PO ca [51] $end
$var wire 1 QO ca [50] $end
$var wire 1 RO ca [49] $end
$var wire 1 SO ca [48] $end
$var wire 1 TO ca [47] $end
$var wire 1 UO ca [46] $end
$var wire 1 VO ca [45] $end
$var wire 1 WO ca [44] $end
$var wire 1 XO ca [43] $end
$var wire 1 YO ca [42] $end
$var wire 1 ZO ca [41] $end
$var wire 1 [O ca [40] $end
$var wire 1 \O ca [39] $end
$var wire 1 ]O ca [38] $end
$var wire 1 ^O ca [37] $end
$var wire 1 _O ca [36] $end
$var wire 1 `O ca [35] $end
$var wire 1 aO ca [34] $end
$var wire 1 bO ca [33] $end
$var wire 1 cO ca [32] $end
$var wire 1 dO ca [31] $end
$var wire 1 eO ca [30] $end
$var wire 1 fO ca [29] $end
$var wire 1 gO ca [28] $end
$var wire 1 hO ca [27] $end
$var wire 1 iO ca [26] $end
$var wire 1 jO ca [25] $end
$var wire 1 kO ca [24] $end
$var wire 1 lO ca [23] $end
$var wire 1 mO ca [22] $end
$var wire 1 nO ca [21] $end
$var wire 1 oO ca [20] $end
$var wire 1 pO ca [19] $end
$var wire 1 qO ca [18] $end
$var wire 1 rO ca [17] $end
$var wire 1 sO ca [16] $end
$var wire 1 tO ca [15] $end
$var wire 1 uO ca [14] $end
$var wire 1 vO ca [13] $end
$var wire 1 wO ca [12] $end
$var wire 1 xO ca [11] $end
$var wire 1 yO ca [10] $end
$var wire 1 zO ca [9] $end
$var wire 1 {O ca [8] $end
$var wire 1 |O ca [7] $end
$var wire 1 }O ca [6] $end
$var wire 1 ~O ca [5] $end
$var wire 1 !P ca [4] $end
$var wire 1 "P ca [3] $end
$var wire 1 #P ca [2] $end
$var wire 1 $P ca [1] $end
$var wire 1 %P ca [0] $end
$upscope $end
$upscope $end

$scope module a0 $end
$var parameter 0 GX BEGINTIME $end
$var wire 1 $ m [63] $end
$var wire 1 % m [62] $end
$var wire 1 & m [61] $end
$var wire 1 ' m [60] $end
$var wire 1 ( m [59] $end
$var wire 1 ) m [58] $end
$var wire 1 * m [57] $end
$var wire 1 + m [56] $end
$var wire 1 , m [55] $end
$var wire 1 - m [54] $end
$var wire 1 . m [53] $end
$var wire 1 / m [52] $end
$var wire 1 0 m [51] $end
$var wire 1 1 m [50] $end
$var wire 1 2 m [49] $end
$var wire 1 3 m [48] $end
$var wire 1 4 m [47] $end
$var wire 1 5 m [46] $end
$var wire 1 6 m [45] $end
$var wire 1 7 m [44] $end
$var wire 1 8 m [43] $end
$var wire 1 9 m [42] $end
$var wire 1 : m [41] $end
$var wire 1 ; m [40] $end
$var wire 1 < m [39] $end
$var wire 1 = m [38] $end
$var wire 1 > m [37] $end
$var wire 1 ? m [36] $end
$var wire 1 @ m [35] $end
$var wire 1 A m [34] $end
$var wire 1 B m [33] $end
$var wire 1 C m [32] $end
$var wire 1 D m [31] $end
$var wire 1 E m [30] $end
$var wire 1 F m [29] $end
$var wire 1 G m [28] $end
$var wire 1 H m [27] $end
$var wire 1 I m [26] $end
$var wire 1 J m [25] $end
$var wire 1 K m [24] $end
$var wire 1 L m [23] $end
$var wire 1 M m [22] $end
$var wire 1 N m [21] $end
$var wire 1 O m [20] $end
$var wire 1 P m [19] $end
$var wire 1 Q m [18] $end
$var wire 1 R m [17] $end
$var wire 1 S m [16] $end
$var wire 1 T m [15] $end
$var wire 1 U m [14] $end
$var wire 1 V m [13] $end
$var wire 1 W m [12] $end
$var wire 1 X m [11] $end
$var wire 1 Y m [10] $end
$var wire 1 Z m [9] $end
$var wire 1 [ m [8] $end
$var wire 1 \ m [7] $end
$var wire 1 ] m [6] $end
$var wire 1 ^ m [5] $end
$var wire 1 _ m [4] $end
$var wire 1 ` m [3] $end
$var wire 1 a m [2] $end
$var wire 1 b m [1] $end
$var wire 1 c m [0] $end
$var wire 1 HX a [31] $end
$var wire 1 IX a [30] $end
$var wire 1 JX a [29] $end
$var wire 1 KX a [28] $end
$var wire 1 LX a [27] $end
$var wire 1 MX a [26] $end
$var wire 1 NX a [25] $end
$var wire 1 OX a [24] $end
$var wire 1 PX a [23] $end
$var wire 1 QX a [22] $end
$var wire 1 RX a [21] $end
$var wire 1 SX a [20] $end
$var wire 1 TX a [19] $end
$var wire 1 UX a [18] $end
$var wire 1 VX a [17] $end
$var wire 1 WX a [16] $end
$var wire 1 XX a [15] $end
$var wire 1 YX a [14] $end
$var wire 1 ZX a [13] $end
$var wire 1 [X a [12] $end
$var wire 1 \X a [11] $end
$var wire 1 ]X a [10] $end
$var wire 1 ^X a [9] $end
$var wire 1 _X a [8] $end
$var wire 1 `X a [7] $end
$var wire 1 aX a [6] $end
$var wire 1 bX a [5] $end
$var wire 1 cX a [4] $end
$var wire 1 dX a [3] $end
$var wire 1 eX a [2] $end
$var wire 1 fX a [1] $end
$var wire 1 gX a [0] $end
$var wire 1 hX b [31] $end
$var wire 1 iX b [30] $end
$var wire 1 jX b [29] $end
$var wire 1 kX b [28] $end
$var wire 1 lX b [27] $end
$var wire 1 mX b [26] $end
$var wire 1 nX b [25] $end
$var wire 1 oX b [24] $end
$var wire 1 pX b [23] $end
$var wire 1 qX b [22] $end
$var wire 1 rX b [21] $end
$var wire 1 sX b [20] $end
$var wire 1 tX b [19] $end
$var wire 1 uX b [18] $end
$var wire 1 vX b [17] $end
$var wire 1 wX b [16] $end
$var wire 1 xX b [15] $end
$var wire 1 yX b [14] $end
$var wire 1 zX b [13] $end
$var wire 1 {X b [12] $end
$var wire 1 |X b [11] $end
$var wire 1 }X b [10] $end
$var wire 1 ~X b [9] $end
$var wire 1 !Y b [8] $end
$var wire 1 "Y b [7] $end
$var wire 1 #Y b [6] $end
$var wire 1 $Y b [5] $end
$var wire 1 %Y b [4] $end
$var wire 1 &Y b [3] $end
$var wire 1 'Y b [2] $end
$var wire 1 (Y b [1] $end
$var wire 1 )Y b [0] $end
$var wire 1 *Y golden_model [63] $end
$var wire 1 +Y golden_model [62] $end
$var wire 1 ,Y golden_model [61] $end
$var wire 1 -Y golden_model [60] $end
$var wire 1 .Y golden_model [59] $end
$var wire 1 /Y golden_model [58] $end
$var wire 1 0Y golden_model [57] $end
$var wire 1 1Y golden_model [56] $end
$var wire 1 2Y golden_model [55] $end
$var wire 1 3Y golden_model [54] $end
$var wire 1 4Y golden_model [53] $end
$var wire 1 5Y golden_model [52] $end
$var wire 1 6Y golden_model [51] $end
$var wire 1 7Y golden_model [50] $end
$var wire 1 8Y golden_model [49] $end
$var wire 1 9Y golden_model [48] $end
$var wire 1 :Y golden_model [47] $end
$var wire 1 ;Y golden_model [46] $end
$var wire 1 <Y golden_model [45] $end
$var wire 1 =Y golden_model [44] $end
$var wire 1 >Y golden_model [43] $end
$var wire 1 ?Y golden_model [42] $end
$var wire 1 @Y golden_model [41] $end
$var wire 1 AY golden_model [40] $end
$var wire 1 BY golden_model [39] $end
$var wire 1 CY golden_model [38] $end
$var wire 1 DY golden_model [37] $end
$var wire 1 EY golden_model [36] $end
$var wire 1 FY golden_model [35] $end
$var wire 1 GY golden_model [34] $end
$var wire 1 HY golden_model [33] $end
$var wire 1 IY golden_model [32] $end
$var wire 1 JY golden_model [31] $end
$var wire 1 KY golden_model [30] $end
$var wire 1 LY golden_model [29] $end
$var wire 1 MY golden_model [28] $end
$var wire 1 NY golden_model [27] $end
$var wire 1 OY golden_model [26] $end
$var wire 1 PY golden_model [25] $end
$var wire 1 QY golden_model [24] $end
$var wire 1 RY golden_model [23] $end
$var wire 1 SY golden_model [22] $end
$var wire 1 TY golden_model [21] $end
$var wire 1 UY golden_model [20] $end
$var wire 1 VY golden_model [19] $end
$var wire 1 WY golden_model [18] $end
$var wire 1 XY golden_model [17] $end
$var wire 1 YY golden_model [16] $end
$var wire 1 ZY golden_model [15] $end
$var wire 1 [Y golden_model [14] $end
$var wire 1 \Y golden_model [13] $end
$var wire 1 ]Y golden_model [12] $end
$var wire 1 ^Y golden_model [11] $end
$var wire 1 _Y golden_model [10] $end
$var wire 1 `Y golden_model [9] $end
$var wire 1 aY golden_model [8] $end
$var wire 1 bY golden_model [7] $end
$var wire 1 cY golden_model [6] $end
$var wire 1 dY golden_model [5] $end
$var wire 1 eY golden_model [4] $end
$var wire 1 fY golden_model [3] $end
$var wire 1 gY golden_model [2] $end
$var wire 1 hY golden_model [1] $end
$var wire 1 iY golden_model [0] $end
$var wire 1 jY test $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0"
1#
b0 d
b0 e
bx H!
bx I!
bx J!
bx K!
bx L!
bx M!
bx N!
bx O!
bx P!
bx Q!
bx R!
bx S!
b0 KQ
b0 LQ
1MQ
b0 NQ
b0 OQ
1PQ
b0 QQ
b0 RQ
1SQ
b0 TQ
b0 UQ
1VQ
b0 WQ
b0 XQ
1YQ
b0 ZQ
b0 [Q
1\Q
b0 ]Q
b0 ^Q
1_Q
b0 `Q
b0 aQ
1bQ
b0 cQ
b0 dQ
1eQ
b0 fQ
b0 gQ
1hQ
b0 iQ
b0 jQ
1kQ
b0 lQ
b0 mQ
1nQ
b0 oQ
b0 pQ
1qQ
b0 rQ
b0 sQ
1tQ
b0 uQ
b0 vQ
1wQ
b0 xQ
b0 yQ
1zQ
bx N:
bx O:
bx P:
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 Q:
bx R:
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 S:
bx T:
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 U:
bx V:
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 W:
bx X:
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 Y:
bx "F
bx0 #F
bx $F
bx0 %F
bx &F
bx0 'F
bx xK
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx0 yK
bx zK
bx00000000000 {K
bx HQ
bx0 IQ
b1111111111111111111111111111111 !
b100100 {Q
b101000 |Q
b101000 }Q
b101000 ~Q
b101000 !R
b100110 "R
b101011 #R
b101111 GS
b101100 wT
b110111 @V
b110111 AV
b1000000 BV
r3.6 GX
xc
xb
xa
x`
x_
x^
x]
x\
x[
xZ
xY
xX
xW
xV
xU
xT
xS
xR
xQ
xP
xO
xN
xM
xL
xK
xJ
xI
xH
xG
xF
xE
xD
xC
xB
xA
x@
x?
x>
x=
x<
x;
x:
x9
x8
x7
x6
x5
x4
x3
x2
x1
x0
x/
x.
x-
x,
x+
x*
x)
x(
x'
x&
x%
x$
0G!
0F!
0E!
0D!
0C!
0B!
0A!
0@!
0?!
0>!
0=!
0<!
0;!
0:!
09!
08!
07!
06!
05!
04!
03!
02!
01!
00!
0/!
0.!
0-!
0,!
0+!
0*!
0)!
0(!
0'!
0&!
0%!
0$!
0#!
0"!
0!!
0~
0}
0|
0{
0z
0y
0x
0w
0v
0u
0t
0s
0r
0q
0p
0o
0n
0m
0l
0k
0j
0i
0h
0g
0f
0X"
0W"
0V"
0U"
0T"
0S"
0R"
0Q"
0P"
0O"
0N"
0M"
0L"
0K"
0J"
0I"
0H"
0G"
0F"
0E"
0D"
0C"
0B"
0A"
0@"
0?"
0>"
0="
0<"
0;"
0:"
09"
08"
0y"
0x"
0w"
0v"
0u"
0t"
0s"
0r"
0q"
0p"
0o"
0n"
0m"
0l"
0k"
0j"
0i"
0h"
0g"
0f"
0e"
0d"
0c"
0b"
0a"
0`"
0_"
0^"
0]"
0\"
0["
0Z"
0Y"
0<#
0;#
0:#
09#
08#
07#
06#
05#
04#
03#
02#
01#
00#
0/#
0.#
0-#
0,#
0+#
0*#
0)#
0(#
0'#
0&#
0%#
0$#
0##
0"#
0!#
0~"
0}"
0|"
0{"
0z"
0]#
0\#
0[#
0Z#
0Y#
0X#
0W#
0V#
0U#
0T#
0S#
0R#
0Q#
0P#
0O#
0N#
0M#
0L#
0K#
0J#
0I#
0H#
0G#
0F#
0E#
0D#
0C#
0B#
0A#
0@#
0?#
0>#
0=#
0~#
0}#
0|#
0{#
0z#
0y#
0x#
0w#
0v#
0u#
0t#
0s#
0r#
0q#
0p#
0o#
0n#
0m#
0l#
0k#
0j#
0i#
0h#
0g#
0f#
0e#
0d#
0c#
0b#
0a#
0`#
0_#
0^#
0A$
0@$
0?$
0>$
0=$
0<$
0;$
0:$
09$
08$
07$
06$
05$
04$
03$
02$
01$
00$
0/$
0.$
0-$
0,$
0+$
0*$
0)$
0($
0'$
0&$
0%$
0$$
0#$
0"$
0!$
0b$
0a$
0`$
0_$
0^$
0]$
0\$
0[$
0Z$
0Y$
0X$
0W$
0V$
0U$
0T$
0S$
0R$
0Q$
0P$
0O$
0N$
0M$
0L$
0K$
0J$
0I$
0H$
0G$
0F$
0E$
0D$
0C$
0B$
0%%
0$%
0#%
0"%
0!%
0~$
0}$
0|$
0{$
0z$
0y$
0x$
0w$
0v$
0u$
0t$
0s$
0r$
0q$
0p$
0o$
0n$
0m$
0l$
0k$
0j$
0i$
0h$
0g$
0f$
0e$
0d$
0c$
0F%
0E%
0D%
0C%
0B%
0A%
0@%
0?%
0>%
0=%
0<%
0;%
0:%
09%
08%
07%
06%
05%
04%
03%
02%
01%
00%
0/%
0.%
0-%
0,%
0+%
0*%
0)%
0(%
0'%
0&%
0g%
0f%
0e%
0d%
0c%
0b%
0a%
0`%
0_%
0^%
0]%
0\%
0[%
0Z%
0Y%
0X%
0W%
0V%
0U%
0T%
0S%
0R%
0Q%
0P%
0O%
0N%
0M%
0L%
0K%
0J%
0I%
0H%
0G%
0*&
0)&
0(&
0'&
0&&
0%&
0$&
0#&
0"&
0!&
0~%
0}%
0|%
0{%
0z%
0y%
0x%
0w%
0v%
0u%
0t%
0s%
0r%
0q%
0p%
0o%
0n%
0m%
0l%
0k%
0j%
0i%
0h%
0K&
0J&
0I&
0H&
0G&
0F&
0E&
0D&
0C&
0B&
0A&
0@&
0?&
0>&
0=&
0<&
0;&
0:&
09&
08&
07&
06&
05&
04&
03&
02&
01&
00&
0/&
0.&
0-&
0,&
0+&
0l&
0k&
0j&
0i&
0h&
0g&
0f&
0e&
0d&
0c&
0b&
0a&
0`&
0_&
0^&
0]&
0\&
0[&
0Z&
0Y&
0X&
0W&
0V&
0U&
0T&
0S&
0R&
0Q&
0P&
0O&
0N&
0M&
0L&
0/'
0.'
0-'
0,'
0+'
0*'
0)'
0('
0''
0&'
0%'
0$'
0#'
0"'
0!'
0~&
0}&
0|&
0{&
0z&
0y&
0x&
0w&
0v&
0u&
0t&
0s&
0r&
0q&
0p&
0o&
0n&
0m&
0P'
0O'
0N'
0M'
0L'
0K'
0J'
0I'
0H'
0G'
0F'
0E'
0D'
0C'
0B'
0A'
0@'
0?'
0>'
0='
0<'
0;'
0:'
09'
08'
07'
06'
05'
04'
03'
02'
01'
00'
0q'
0p'
0o'
0n'
0m'
0l'
0k'
0j'
0i'
0h'
0g'
0f'
0e'
0d'
0c'
0b'
0a'
0`'
0_'
0^'
0]'
0\'
0['
0Z'
0Y'
0X'
0W'
0V'
0U'
0T'
0S'
0R'
0Q'
02(
01(
00(
0/(
0.(
0-(
0,(
0+(
0*(
0)(
0((
0'(
0&(
0%(
0$(
0#(
0"(
0!(
0~'
0}'
0|'
0{'
0z'
0y'
0x'
0w'
0v'
0u'
0t'
0s'
0r'
04(
03(
06(
05(
08(
07(
0:(
09(
0<(
0;(
0>(
0=(
0@(
0?(
0B(
0A(
0D(
0C(
0F(
0E(
0H(
0G(
0J(
0I(
0L(
0K(
0N(
0M(
0P(
0O(
0R(
0Q(
0r(
0q(
0p(
0o(
0n(
0m(
0l(
0k(
0j(
0i(
0h(
0g(
0f(
0e(
0d(
0c(
0b(
0a(
0`(
0_(
0^(
0](
0\(
0[(
0Z(
0Y(
0X(
0W(
0V(
0U(
0T(
0S(
1%)
1$)
1#)
1")
1!)
1~(
1}(
1|(
1{(
1z(
1y(
1x(
1w(
1v(
1u(
1t(
zs(
0I)
0H)
0G)
0F)
0E)
0D)
0C)
0B)
0A)
0@)
0?)
0>)
0=)
0<)
0;)
0:)
09)
08)
07)
06)
05)
04)
03)
02)
01)
00)
0/)
0.)
0-)
0,)
0+)
0*)
0))
0()
0')
0&)
0m)
0l)
0k)
0j)
0i)
0h)
0g)
0f)
0e)
0d)
0c)
0b)
0a)
0`)
0_)
0^)
0])
0\)
0[)
0Z)
0Y)
0X)
0W)
0V)
0U)
0T)
0S)
0R)
0Q)
0P)
0O)
0N)
0M)
0L)
0K)
1J)
03*
02*
01*
00*
0/*
0.*
0-*
0,*
0+*
0**
0)*
0(*
0'*
0&*
0%*
0$*
0#*
0"*
0!*
0~)
0})
0|)
0{)
0z)
0y)
0x)
0w)
0v)
0u)
0t)
0s)
0r)
0q)
0p)
0o)
1n)
zW*
zV*
zU*
zT*
zS*
zR*
zQ*
zP*
zO*
zN*
zM*
zL*
zK*
zJ*
zI*
zH*
zG*
zF*
zE*
zD*
zC*
zB*
zA*
z@*
z?*
z>*
z=*
z<*
z;*
z:*
z9*
z8*
z7*
z6*
z5*
z4*
z{*
zz*
zy*
zx*
zw*
zv*
zu*
zt*
zs*
zr*
zq*
zp*
zo*
zn*
zm*
zl*
zk*
zj*
zi*
zh*
zg*
zf*
ze*
zd*
zc*
zb*
za*
z`*
z_*
z^*
z]*
z\*
z[*
zZ*
zY*
zX*
0A+
0@+
0?+
0>+
0=+
0<+
0;+
0:+
09+
08+
07+
06+
05+
04+
03+
02+
01+
00+
0/+
0.+
0-+
0,+
0++
0*+
0)+
0(+
0'+
0&+
0%+
0$+
0#+
0"+
0!+
0~*
0}*
0|*
0e+
0d+
0c+
0b+
0a+
0`+
0_+
0^+
0]+
0\+
0[+
0Z+
0Y+
0X+
0W+
0V+
0U+
0T+
0S+
0R+
0Q+
0P+
0O+
0N+
0M+
0L+
0K+
0J+
0I+
0H+
0G+
0F+
0E+
0D+
0C+
1B+
0/,
0.,
0-,
0,,
0+,
0*,
0),
0(,
0',
0&,
0%,
0$,
0#,
0",
0!,
0~+
0}+
0|+
0{+
0z+
0y+
0x+
0w+
0v+
0u+
0t+
0s+
0r+
0q+
0p+
0o+
0n+
0m+
0l+
0k+
1j+
0i+
0h+
0g+
0f+
0W,
0V,
0U,
0T,
0S,
0R,
0Q,
0P,
0O,
0N,
0M,
0L,
0K,
0J,
0I,
0H,
0G,
0F,
0E,
0D,
0C,
0B,
0A,
0@,
0?,
0>,
0=,
0<,
0;,
0:,
09,
08,
07,
06,
05,
04,
03,
12,
01,
00,
0!-
0~,
0},
0|,
0{,
0z,
0y,
0x,
0w,
0v,
0u,
0t,
0s,
0r,
0q,
0p,
0o,
0n,
0m,
0l,
0k,
0j,
0i,
0h,
0g,
0f,
0e,
0d,
0c,
0b,
0a,
0`,
0_,
0^,
0],
0\,
0[,
0Z,
0Y,
1X,
zI-
zH-
zG-
zF-
zE-
zD-
zC-
zB-
zA-
z@-
z?-
z>-
z=-
z<-
z;-
z:-
z9-
z8-
z7-
z6-
z5-
z4-
z3-
z2-
z1-
z0-
z/-
z.-
z--
z,-
z+-
z*-
z)-
z(-
z'-
z&-
z%-
z$-
z#-
z"-
zq-
zp-
zo-
zn-
zm-
zl-
zk-
zj-
zi-
zh-
zg-
zf-
ze-
zd-
zc-
zb-
za-
z`-
z_-
z^-
z]-
z\-
z[-
zZ-
zY-
zX-
zW-
zV-
zU-
zT-
zS-
zR-
zQ-
zP-
zO-
zN-
zM-
zL-
zK-
zJ-
0;.
0:.
09.
08.
07.
06.
05.
04.
03.
02.
01.
00.
0/.
0..
0-.
0,.
0+.
0*.
0).
0(.
0'.
0&.
0%.
0$.
0#.
0".
0!.
0~-
0}-
0|-
0{-
0z-
0y-
0x-
0w-
1v-
0u-
1t-
0s-
1r-
0c.
0b.
0a.
0`.
0_.
0^.
0].
0\.
0[.
0Z.
0Y.
0X.
0W.
0V.
0U.
0T.
0S.
0R.
0Q.
0P.
0O.
0N.
0M.
0L.
0K.
0J.
0I.
0H.
0G.
0F.
0E.
0D.
0C.
0B.
0A.
0@.
0?.
0>.
0=.
0<.
0-/
0,/
0+/
0*/
0)/
0(/
0'/
0&/
0%/
0$/
0#/
0"/
0!/
0~.
0}.
0|.
0{.
0z.
0y.
0x.
0w.
0v.
0u.
0t.
0s.
0r.
0q.
0p.
0o.
0n.
0m.
0l.
0k.
0j.
0i.
1h.
0g.
0f.
0e.
0d.
0U/
0T/
0S/
0R/
0Q/
0P/
0O/
0N/
0M/
0L/
0K/
0J/
0I/
0H/
0G/
0F/
0E/
0D/
0C/
0B/
0A/
0@/
0?/
0>/
0=/
0</
0;/
0:/
09/
08/
07/
06/
05/
04/
03/
02/
01/
10/
0//
0./
0}/
0|/
0{/
0z/
0y/
0x/
0w/
0v/
0u/
0t/
0s/
0r/
0q/
0p/
0o/
0n/
0m/
0l/
0k/
0j/
0i/
0h/
0g/
0f/
0e/
0d/
0c/
0b/
0a/
0`/
0_/
0^/
0]/
0\/
0[/
0Z/
0Y/
0X/
0W/
1V/
zG0
zF0
zE0
zD0
zC0
zB0
zA0
z@0
z?0
z>0
z=0
z<0
z;0
z:0
z90
z80
z70
z60
z50
z40
z30
z20
z10
z00
z/0
z.0
z-0
z,0
z+0
z*0
z)0
z(0
z'0
z&0
z%0
z$0
z#0
z"0
z!0
z~/
zo0
zn0
zm0
zl0
zk0
zj0
zi0
zh0
zg0
zf0
ze0
zd0
zc0
zb0
za0
z`0
z_0
z^0
z]0
z\0
z[0
zZ0
zY0
zX0
zW0
zV0
zU0
zT0
zS0
zR0
zQ0
zP0
zO0
zN0
zM0
zL0
zK0
zJ0
zI0
zH0
091
081
071
061
051
041
031
021
011
001
0/1
0.1
0-1
0,1
0+1
0*1
0)1
0(1
0'1
0&1
0%1
0$1
0#1
0"1
0!1
0~0
0}0
0|0
0{0
0z0
0y0
0x0
0w0
0v0
0u0
1t0
0s0
1r0
0q0
1p0
0a1
0`1
0_1
0^1
0]1
0\1
0[1
0Z1
0Y1
0X1
0W1
0V1
0U1
0T1
0S1
0R1
0Q1
0P1
0O1
0N1
0M1
0L1
0K1
0J1
0I1
0H1
0G1
0F1
0E1
0D1
0C1
0B1
0A1
0@1
0?1
0>1
0=1
0<1
0;1
0:1
0+2
0*2
0)2
0(2
0'2
0&2
0%2
0$2
0#2
0"2
0!2
0~1
0}1
0|1
0{1
0z1
0y1
0x1
0w1
0v1
0u1
0t1
0s1
0r1
0q1
0p1
0o1
0n1
0m1
0l1
0k1
0j1
0i1
0h1
0g1
1f1
0e1
0d1
0c1
0b1
0S2
0R2
0Q2
0P2
0O2
0N2
0M2
0L2
0K2
0J2
0I2
0H2
0G2
0F2
0E2
0D2
0C2
0B2
0A2
0@2
0?2
0>2
0=2
0<2
0;2
0:2
092
082
072
062
052
042
032
022
012
002
0/2
1.2
0-2
0,2
0{2
0z2
0y2
0x2
0w2
0v2
0u2
0t2
0s2
0r2
0q2
0p2
0o2
0n2
0m2
0l2
0k2
0j2
0i2
0h2
0g2
0f2
0e2
0d2
0c2
0b2
0a2
0`2
0_2
0^2
0]2
0\2
0[2
0Z2
0Y2
0X2
0W2
0V2
0U2
1T2
zE3
zD3
zC3
zB3
zA3
z@3
z?3
z>3
z=3
z<3
z;3
z:3
z93
z83
z73
z63
z53
z43
z33
z23
z13
z03
z/3
z.3
z-3
z,3
z+3
z*3
z)3
z(3
z'3
z&3
z%3
z$3
z#3
z"3
z!3
z~2
z}2
z|2
zm3
zl3
zk3
zj3
zi3
zh3
zg3
zf3
ze3
zd3
zc3
zb3
za3
z`3
z_3
z^3
z]3
z\3
z[3
zZ3
zY3
zX3
zW3
zV3
zU3
zT3
zS3
zR3
zQ3
zP3
zO3
zN3
zM3
zL3
zK3
zJ3
zI3
zH3
zG3
zF3
074
064
054
044
034
024
014
004
0/4
0.4
0-4
0,4
0+4
0*4
0)4
0(4
0'4
0&4
0%4
0$4
0#4
0"4
0!4
0~3
0}3
0|3
0{3
0z3
0y3
0x3
0w3
0v3
0u3
0t3
0s3
1r3
0q3
1p3
0o3
1n3
0_4
0^4
0]4
0\4
0[4
0Z4
0Y4
0X4
0W4
0V4
0U4
0T4
0S4
0R4
0Q4
0P4
0O4
0N4
0M4
0L4
0K4
0J4
0I4
0H4
0G4
0F4
0E4
0D4
0C4
0B4
0A4
0@4
0?4
0>4
0=4
0<4
0;4
0:4
094
084
0)5
0(5
0'5
0&5
0%5
0$5
0#5
0"5
0!5
0~4
0}4
0|4
0{4
0z4
0y4
0x4
0w4
0v4
0u4
0t4
0s4
0r4
0q4
0p4
0o4
0n4
0m4
0l4
0k4
0j4
0i4
0h4
0g4
0f4
0e4
1d4
0c4
0b4
0a4
0`4
0Q5
0P5
0O5
0N5
0M5
0L5
0K5
0J5
0I5
0H5
0G5
0F5
0E5
0D5
0C5
0B5
0A5
0@5
0?5
0>5
0=5
0<5
0;5
0:5
095
085
075
065
055
045
035
025
015
005
0/5
0.5
0-5
1,5
0+5
0*5
0y5
0x5
0w5
0v5
0u5
0t5
0s5
0r5
0q5
0p5
0o5
0n5
0m5
0l5
0k5
0j5
0i5
0h5
0g5
0f5
0e5
0d5
0c5
0b5
0a5
0`5
0_5
0^5
0]5
0\5
0[5
0Z5
0Y5
0X5
0W5
0V5
0U5
0T5
0S5
1R5
zC6
zB6
zA6
z@6
z?6
z>6
z=6
z<6
z;6
z:6
z96
z86
z76
z66
z56
z46
z36
z26
z16
z06
z/6
z.6
z-6
z,6
z+6
z*6
z)6
z(6
z'6
z&6
z%6
z$6
z#6
z"6
z!6
z~5
z}5
z|5
z{5
zz5
zk6
zj6
zi6
zh6
zg6
zf6
ze6
zd6
zc6
zb6
za6
z`6
z_6
z^6
z]6
z\6
z[6
zZ6
zY6
zX6
zW6
zV6
zU6
zT6
zS6
zR6
zQ6
zP6
zO6
zN6
zM6
zL6
zK6
zJ6
zI6
zH6
zG6
zF6
zE6
zD6
057
047
037
027
017
007
0/7
0.7
0-7
0,7
0+7
0*7
0)7
0(7
0'7
0&7
0%7
0$7
0#7
0"7
0!7
0~6
0}6
0|6
0{6
0z6
0y6
0x6
0w6
0v6
0u6
0t6
0s6
0r6
0q6
1p6
0o6
1n6
0m6
1l6
0]7
0\7
0[7
0Z7
0Y7
0X7
0W7
0V7
0U7
0T7
0S7
0R7
0Q7
0P7
0O7
0N7
0M7
0L7
0K7
0J7
0I7
0H7
0G7
0F7
0E7
0D7
0C7
0B7
0A7
0@7
0?7
0>7
0=7
0<7
0;7
0:7
097
087
077
067
0%8
0$8
0#8
0"8
0!8
0~7
0}7
0|7
0{7
0z7
0y7
0x7
0w7
0v7
0u7
0t7
0s7
0r7
0q7
0p7
0o7
0n7
0m7
0l7
0k7
0j7
0i7
0h7
0g7
0f7
0e7
0d7
0c7
0b7
0a7
1`7
0_7
0^7
0K8
0J8
0I8
0H8
0G8
0F8
0E8
0D8
0C8
0B8
0A8
0@8
0?8
0>8
0=8
0<8
0;8
0:8
098
088
078
068
058
048
038
028
018
008
0/8
0.8
0-8
0,8
0+8
0*8
0)8
0(8
0'8
1&8
0q8
0p8
0o8
0n8
0m8
0l8
0k8
0j8
0i8
0h8
1g8
0f8
1e8
0d8
1c8
0b8
1a8
0`8
1_8
0^8
1]8
0\8
1[8
0Z8
1Y8
0X8
1W8
0V8
1U8
0T8
1S8
0R8
1Q8
0P8
1O8
0N8
1M8
0L8
z99
z89
z79
z69
z59
z49
z39
z29
z19
z09
z/9
z.9
z-9
z,9
z+9
z*9
z)9
z(9
z'9
z&9
z%9
z$9
z#9
z"9
z!9
z~8
z}8
z|8
z{8
zz8
zy8
zx8
zw8
zv8
zu8
zt8
zs8
zr8
z_9
z^9
z]9
z\9
z[9
zZ9
zY9
zX9
zW9
zV9
zU9
zT9
zS9
zR9
zQ9
zP9
zO9
zN9
zM9
zL9
zK9
zJ9
zI9
zH9
zG9
zF9
zE9
zD9
zC9
zB9
zA9
z@9
z?9
z>9
z=9
z<9
z;9
z:9
0':
0&:
0%:
0$:
0#:
0":
0!:
0~9
0}9
0|9
1{9
0z9
1y9
0x9
1w9
0v9
1u9
0t9
1s9
0r9
1q9
0p9
1o9
0n9
1m9
0l9
1k9
0j9
1i9
0h9
1g9
0f9
1e9
0d9
1c9
1b9
1a9
1`9
0M:
0L:
0K:
0J:
0I:
0H:
0G:
0F:
0E:
0D:
0C:
0B:
0A:
0@:
0?:
0>:
0=:
0<:
0;:
0::
09:
08:
07:
06:
05:
04:
03:
02:
01:
00:
0/:
0.:
0-:
0,:
0+:
0*:
0):
0(:
x&;
x%;
x$;
x#;
x";
x!;
x~:
x}:
x|:
x{:
xz:
xy:
xx:
xw:
xv:
xu:
xt:
xs:
xr:
xq:
xp:
xo:
xn:
xm:
xl:
xk:
xj:
xi:
xh:
xg:
xf:
xe:
xd:
xc:
xb:
xa:
0`:
0_:
0^:
0]:
0\:
0[:
0Z:
0Q;
xP;
xO;
xN;
xM;
xL;
xK;
xJ;
xI;
xH;
xG;
xF;
xE;
xD;
xC;
xB;
xA;
x@;
x?;
x>;
x=;
x<;
x;;
x:;
x9;
x8;
x7;
x6;
x5;
x4;
x3;
x2;
x1;
x0;
x/;
x.;
x-;
0,;
0+;
0*;
0);
0(;
0';
0|;
0{;
xz;
xy;
xx;
xw;
xv;
xu;
xt;
xs;
xr;
xq;
xp;
xo;
xn;
xm;
xl;
xk;
xj;
xi;
xh;
xg;
xf;
xe;
xd;
xc;
xb;
xa;
x`;
x_;
x^;
x];
x\;
x[;
xZ;
xY;
xX;
xW;
xV;
xU;
xT;
xS;
0R;
0I<
0H<
0G<
0F<
0E<
xD<
xC<
xB<
xA<
x@<
x?<
x><
x=<
x<<
x;<
x:<
x9<
x8<
x7<
x6<
x5<
x4<
x3<
x2<
x1<
x0<
x/<
x.<
x-<
x,<
x+<
x*<
x)<
x(<
x'<
x&<
x%<
x$<
x#<
x"<
x!<
0~;
0};
0t<
xs<
xr<
xq<
xp<
xo<
xn<
xm<
xl<
xk<
xj<
xi<
xh<
xg<
xf<
xe<
xd<
xc<
xb<
xa<
x`<
x_<
x^<
x]<
x\<
x[<
xZ<
xY<
xX<
xW<
xV<
xU<
xT<
xS<
xR<
xQ<
xP<
xO<
0N<
0M<
0L<
0K<
0J<
xA=
x@=
x?=
x>=
x==
x<=
x;=
x:=
x9=
x8=
x7=
x6=
x5=
x4=
x3=
x2=
x1=
x0=
x/=
x.=
x-=
x,=
x+=
x*=
x)=
x(=
x'=
x&=
x%=
x$=
x#=
x"=
x!=
x~<
x}<
x|<
x{<
0z<
0y<
0x<
0w<
0v<
0u<
xl=
xk=
xj=
xi=
xh=
xg=
xf=
xe=
xd=
xc=
xb=
xa=
x`=
x_=
x^=
x]=
x\=
x[=
xZ=
xY=
xX=
xW=
xV=
xU=
xT=
xS=
xR=
xQ=
xP=
xO=
xN=
xM=
xL=
xK=
xJ=
xI=
xH=
xG=
xF=
xE=
xD=
xC=
0B=
09>
x8>
x7>
x6>
x5>
x4>
x3>
x2>
x1>
x0>
x/>
x.>
x->
x,>
x+>
x*>
x)>
x(>
x'>
x&>
x%>
x$>
x#>
x">
x!>
x~=
x}=
x|=
x{=
xz=
xy=
xx=
xw=
xv=
xu=
xt=
xs=
xr=
xq=
xp=
xo=
0n=
0m=
xh>
xg>
xf>
xe>
xd>
xc>
xb>
xa>
x`>
x_>
x^>
x]>
x\>
x[>
xZ>
xY>
xX>
xW>
xV>
xU>
xT>
xS>
xR>
xQ>
xP>
xO>
xN>
xM>
xL>
xK>
xJ>
xI>
xH>
xG>
xF>
xE>
xD>
xC>
xB>
xA>
0@>
0?>
0>>
0=>
0<>
0;>
0:>
09?
08?
07?
x6?
x5?
x4?
x3?
x2?
x1?
x0?
x/?
x.?
x-?
x,?
x+?
x*?
x)?
x(?
x'?
x&?
x%?
x$?
x#?
x"?
x!?
x~>
x}>
x|>
x{>
xz>
xy>
xx>
xw>
xv>
xu>
xt>
xs>
xr>
xq>
0p>
0o>
0n>
0m>
0l>
0k>
0j>
0i>
0h?
0g?
0f?
0e?
0d?
0c?
xb?
xa?
x`?
x_?
x^?
x]?
x\?
x[?
xZ?
xY?
xX?
xW?
xV?
xU?
xT?
xS?
xR?
xQ?
xP?
xO?
xN?
xM?
xL?
xK?
xJ?
xI?
xH?
xG?
xF?
xE?
xD?
xC?
xB?
xA?
x@?
x??
x>?
x=?
x<?
x;?
0:?
09@
08@
07@
06@
05@
04@
03@
02@
01@
x0@
x/@
x.@
x-@
x,@
x+@
x*@
x)@
x(@
x'@
x&@
x%@
x$@
x#@
x"@
x!@
x~?
x}?
x|?
x{?
xz?
xy?
xx?
xw?
xv?
xu?
xt?
xs?
xr?
xq?
xp?
xo?
xn?
xm?
xl?
xk?
0j?
0i?
0h@
xg@
xf@
xe@
xd@
xc@
xb@
xa@
x`@
x_@
x^@
x]@
x\@
x[@
xZ@
xY@
xX@
xW@
xV@
xU@
xT@
xS@
xR@
xQ@
xP@
xO@
xN@
xM@
xL@
xK@
xJ@
xI@
xH@
xG@
xF@
xE@
xD@
xC@
xB@
xA@
x@@
0?@
0>@
0=@
0<@
0;@
0:@
x9A
x8A
x7A
x6A
x5A
x4A
x3A
x2A
x1A
x0A
x/A
x.A
x-A
x,A
x+A
x*A
x)A
x(A
x'A
x&A
x%A
x$A
x#A
x"A
x!A
x~@
x}@
x|@
x{@
xz@
xy@
xx@
xw@
xv@
xu@
xt@
xs@
xr@
xq@
xp@
0o@
0n@
0m@
0l@
0k@
0j@
0i@
xhA
xgA
xfA
xeA
xdA
xcA
xbA
xaA
x`A
x_A
x^A
x]A
x\A
x[A
xZA
xYA
xXA
xWA
xVA
xUA
xTA
xSA
xRA
xQA
xPA
xOA
xNA
xMA
xLA
xKA
xJA
xIA
xHA
xGA
xFA
xEA
xDA
xCA
xBA
xAA
x@A
x?A
x>A
x=A
x<A
x;A
0:A
09B
x8B
x7B
x6B
x5B
x4B
x3B
x2B
x1B
x0B
x/B
x.B
x-B
x,B
x+B
x*B
x)B
x(B
x'B
x&B
x%B
x$B
x#B
x"B
x!B
x~A
x}A
x|A
x{A
xzA
xyA
xxA
xwA
xvA
xuA
xtA
xsA
xrA
xqA
xpA
xoA
xnA
xmA
xlA
xkA
0jA
0iA
xeB
xdB
xcB
xbB
xaB
x`B
x_B
x^B
x]B
x\B
x[B
xZB
xYB
xXB
xWB
xVB
xUB
xTB
xSB
xRB
xQB
xPB
xOB
xNB
xMB
xLB
xKB
xJB
xIB
xHB
xGB
xFB
xEB
xDB
xCB
xBB
xAB
x@B
x?B
x>B
0=B
0<B
0;B
0:B
03C
02C
01C
x0C
x/C
x.C
x-C
x,C
x+C
x*C
x)C
x(C
x'C
x&C
x%C
x$C
x#C
x"C
x!C
x~B
x}B
x|B
x{B
xzB
xyB
xxB
xwB
xvB
xuB
xtB
xsB
xrB
xqB
xpB
xoB
xnB
xmB
xlB
xkB
0jB
0iB
0hB
0gB
0fB
0_C
0^C
0]C
0\C
0[C
0ZC
xYC
xXC
xWC
xVC
xUC
xTC
xSC
xRC
xQC
xPC
xOC
xNC
xMC
xLC
xKC
xJC
xIC
xHC
xGC
xFC
xEC
xDC
xCC
xBC
xAC
x@C
x?C
x>C
x=C
x<C
x;C
x:C
x9C
x8C
x7C
x6C
x5C
x4C
0-D
0,D
0+D
0*D
0)D
0(D
0'D
0&D
0%D
x$D
x#D
x"D
x!D
x~C
x}C
x|C
x{C
xzC
xyC
xxC
xwC
xvC
xuC
xtC
xsC
xrC
xqC
xpC
xoC
xnC
xmC
xlC
xkC
xjC
xiC
xhC
xgC
xfC
xeC
xdC
xcC
xbC
xaC
x`C
0YD
xXD
xWD
xVD
xUD
xTD
xSD
xRD
xQD
xPD
xOD
xND
xMD
xLD
xKD
xJD
xID
xHD
xGD
xFD
xED
xDD
xCD
xBD
xAD
x@D
x?D
x>D
x=D
x<D
x;D
x:D
x9D
x8D
x7D
x6D
x5D
x4D
x3D
x2D
x1D
00D
0/D
0.D
x'E
x&E
x%E
x$E
x#E
x"E
x!E
x~D
x}D
x|D
x{D
xzD
xyD
xxD
xwD
xvD
xuD
xtD
xsD
xrD
xqD
xpD
xoD
xnD
xmD
xlD
xkD
xjD
xiD
xhD
xgD
xfD
xeD
xdD
xcD
xbD
xaD
x`D
x_D
x^D
0]D
0\D
0[D
0ZD
xSE
xRE
xQE
xPE
xOE
xNE
xME
xLE
xKE
xJE
xIE
xHE
xGE
xFE
xEE
xDE
xCE
xBE
xAE
x@E
x?E
x>E
x=E
x<E
x;E
x:E
x9E
x8E
x7E
x6E
x5E
x4E
x3E
x2E
x1E
x0E
x/E
x.E
x-E
x,E
x+E
x*E
x)E
x(E
0!F
x~E
x}E
x|E
x{E
xzE
xyE
xxE
xwE
xvE
xuE
xtE
xsE
xrE
xqE
xpE
xoE
xnE
xmE
xlE
xkE
xjE
xiE
xhE
xgE
xfE
xeE
xdE
xcE
xbE
xaE
x`E
x_E
x^E
x]E
x\E
x[E
xZE
xYE
xXE
xWE
xVE
xUE
xTE
xNR
xMR
xLR
xKR
xJR
xIR
xHR
xGR
xFR
xER
xDR
xCR
xBR
xAR
x@R
x?R
x>R
x=R
x<R
x;R
x:R
x9R
x8R
x7R
x6R
x5R
x4R
x3R
x2R
x1R
x0R
x/R
x.R
x-R
x,R
x+R
x*R
0)R
0(R
0'R
0&R
0%R
0$R
0yR
0xR
xwR
xvR
xuR
xtR
xsR
xrR
xqR
xpR
xoR
xnR
xmR
xlR
xkR
xjR
xiR
xhR
xgR
xfR
xeR
xdR
xcR
xbR
xaR
x`R
x_R
x^R
x]R
x\R
x[R
xZR
xYR
xXR
xWR
xVR
xUR
xTR
xSR
xRR
xQR
xPR
0OR
xFS
xES
xDS
xCS
xBS
xAS
x@S
x?S
x>S
x=S
x<S
x;S
x:S
x9S
x8S
x7S
x6S
x5S
x4S
x3S
x2S
x1S
x0S
x/S
x.S
x-S
x,S
x+S
x*S
x)S
x(S
x'S
x&S
x%S
x$S
x#S
x"S
x!S
x~R
x}R
x|R
x{R
0zR
xvS
xuS
xtS
xsS
xrS
xqS
xpS
xoS
xnS
xmS
xlS
xkS
xjS
xiS
xhS
xgS
xfS
xeS
xdS
xcS
xbS
xaS
x`S
x_S
x^S
x]S
x\S
x[S
xZS
xYS
xXS
xWS
xVS
xUS
xTS
xSS
xRS
xQS
xPS
xOS
0NS
0MS
0LS
0KS
0JS
0IS
0HS
0GT
0FT
0ET
0DT
0CT
0BT
xAT
x@T
x?T
x>T
x=T
x<T
x;T
x:T
x9T
x8T
x7T
x6T
x5T
x4T
x3T
x2T
x1T
x0T
x/T
x.T
x-T
x,T
x+T
x*T
x)T
x(T
x'T
x&T
x%T
x$T
x#T
x"T
x!T
x~S
x}S
x|S
x{S
xzS
xyS
xxS
0wS
xvT
xuT
xtT
xsT
xrT
xqT
xpT
xoT
xnT
xmT
xlT
xkT
xjT
xiT
xhT
xgT
xfT
xeT
xdT
xcT
xbT
xaT
x`T
x_T
x^T
x]T
x\T
x[T
xZT
xYT
xXT
xWT
xVT
xUT
xTT
xST
xRT
xQT
xPT
xOT
xNT
xMT
xLT
xKT
xJT
xIT
0HT
xEU
xDU
xCU
xBU
xAU
x@U
x?U
x>U
x=U
x<U
x;U
x:U
x9U
x8U
x7U
x6U
x5U
x4U
x3U
x2U
x1U
x0U
x/U
x.U
x-U
x,U
x+U
x*U
x)U
x(U
x'U
x&U
x%U
x$U
x#U
x"U
x!U
x~T
x}T
x|T
0{T
0zT
0yT
0xT
0qU
0pU
0oU
0nU
0mU
0lU
xkU
xjU
xiU
xhU
xgU
xfU
xeU
xdU
xcU
xbU
xaU
x`U
x_U
x^U
x]U
x\U
x[U
xZU
xYU
xXU
xWU
xVU
xUU
xTU
xSU
xRU
xQU
xPU
xOU
xNU
xMU
xLU
xKU
xJU
xIU
xHU
xGU
xFU
x?V
x>V
x=V
x<V
x;V
x:V
x9V
x8V
x7V
x6V
x5V
x4V
x3V
x2V
x1V
x0V
x/V
x.V
x-V
x,V
x+V
x*V
x)V
x(V
x'V
x&V
x%V
x$V
x#V
x"V
x!V
x~U
x}U
x|U
x{U
xzU
xyU
xxU
xwU
xvU
xuU
xtU
xsU
xrU
x^F
x]F
x\F
x[F
xZF
xYF
xXF
xWF
xVF
xUF
xTF
xSF
xRF
xQF
xPF
xOF
xNF
xMF
xLF
xKF
xJF
xIF
xHF
xGF
xFF
xEF
xDF
xCF
xBF
xAF
x@F
x?F
x>F
x=F
x<F
x;F
x:F
x9F
x8F
x7F
x6F
x5F
x4F
03F
02F
01F
00F
0/F
0.F
0-F
0,F
0+F
0*F
0)F
0(F
07G
06G
x5G
x4G
x3G
x2G
x1G
x0G
x/G
x.G
x-G
x,G
x+G
x*G
x)G
x(G
x'G
x&G
x%G
x$G
x#G
x"G
x!G
x~F
x}F
x|F
x{F
xzF
xyF
xxF
xwF
xvF
xuF
xtF
xsF
xrF
xqF
xpF
xoF
xnF
xmF
xlF
xkF
xjF
0iF
0hF
0gF
0fF
0eF
0dF
0cF
0bF
0aF
0`F
0_F
0nG
0mG
0lG
0kG
0jG
0iG
0hG
0gG
xfG
xeG
xdG
xcG
xbG
xaG
x`G
x_G
x^G
x]G
x\G
x[G
xZG
xYG
xXG
xWG
xVG
xUG
xTG
xSG
xRG
xQG
xPG
xOG
xNG
xMG
xLG
xKG
xJG
xIG
xHG
xGG
xFG
xEG
xDG
xCG
xBG
xAG
x@G
x?G
x>G
x=G
x<G
x;G
x:G
x9G
x8G
xGH
xFH
xEH
xDH
xCH
xBH
xAH
x@H
x?H
x>H
x=H
x<H
x;H
x:H
x9H
x8H
x7H
x6H
x5H
x4H
x3H
x2H
x1H
x0H
x/H
x.H
x-H
x,H
x+H
x*H
x)H
x(H
x'H
x&H
x%H
x$H
x#H
x"H
x!H
x~G
x}G
x|G
x{G
xzG
xyG
xxG
xwG
xvG
xuG
xtG
xsG
xrG
xqG
xpG
xoG
0~H
0}H
x|H
x{H
xzH
xyH
xxH
xwH
xvH
xuH
xtH
xsH
xrH
xqH
xpH
xoH
xnH
xmH
xlH
xkH
xjH
xiH
xhH
xgH
xfH
xeH
xdH
xcH
xbH
xaH
x`H
x_H
x^H
x]H
x\H
x[H
xZH
xYH
xXH
xWH
xVH
xUH
xTH
xSH
0RH
0QH
0PH
0OH
0NH
0MH
0LH
0KH
0JH
0IH
0HH
0WI
xVI
xUI
xTI
xSI
xRI
xQI
xPI
xOI
xNI
xMI
xLI
xKI
xJI
xII
xHI
xGI
xFI
xEI
xDI
xCI
xBI
xAI
x@I
x?I
x>I
x=I
x<I
x;I
x:I
x9I
x8I
x7I
x6I
x5I
x4I
x3I
x2I
x1I
x0I
x/I
x.I
x-I
x,I
x+I
x*I
x)I
0(I
0'I
0&I
0%I
0$I
0#I
0"I
0!I
00J
0/J
0.J
0-J
0,J
0+J
0*J
0)J
0(J
0'J
0&J
x%J
x$J
x#J
x"J
x!J
x~I
x}I
x|I
x{I
xzI
xyI
xxI
xwI
xvI
xuI
xtI
xsI
xrI
xqI
xpI
xoI
xnI
xmI
xlI
xkI
xjI
xiI
xhI
xgI
xfI
xeI
xdI
xcI
xbI
xaI
x`I
x_I
x^I
x]I
x\I
x[I
xZI
xYI
xXI
0gJ
0fJ
0eJ
0dJ
0cJ
0bJ
0aJ
0`J
0_J
0^J
0]J
0\J
0[J
xZJ
xYJ
xXJ
xWJ
xVJ
xUJ
xTJ
xSJ
xRJ
xQJ
xPJ
xOJ
xNJ
xMJ
xLJ
xKJ
xJJ
xIJ
xHJ
xGJ
xFJ
xEJ
xDJ
xCJ
xBJ
xAJ
x@J
x?J
x>J
x=J
x<J
x;J
x:J
x9J
x8J
x7J
x6J
x5J
x4J
x3J
x2J
x1J
0@K
x?K
x>K
x=K
x<K
x;K
x:K
x9K
x8K
x7K
x6K
x5K
x4K
x3K
x2K
x1K
x0K
x/K
x.K
x-K
x,K
x+K
x*K
x)K
x(K
x'K
x&K
x%K
x$K
x#K
x"K
x!K
x~J
x}J
x|J
x{J
xzJ
xyJ
xxJ
xwJ
xvJ
xuJ
xtJ
xsJ
xrJ
xqJ
xpJ
xoJ
xnJ
xmJ
xlJ
xkJ
xjJ
xiJ
xhJ
0wK
0vK
0uK
0tK
0sK
0rK
0qK
0pK
0oK
0nK
0mK
xlK
xkK
xjK
xiK
xhK
xgK
xfK
xeK
xdK
xcK
xbK
xaK
x`K
x_K
x^K
x]K
x\K
x[K
xZK
xYK
xXK
xWK
xVK
xUK
xTK
xSK
xRK
xQK
xPK
xOK
xNK
xMK
xLK
xKK
xJK
xIK
xHK
xGK
xFK
xEK
xDK
xCK
xBK
xAK
x]L
x\L
x[L
xZL
xYL
xXL
xWL
xVL
xUL
xTL
xSL
xRL
xQL
xPL
xOL
xNL
xML
xLL
xKL
xJL
xIL
xHL
xGL
xFL
xEL
xDL
xCL
xBL
xAL
x@L
x?L
x>L
x=L
x<L
x;L
x:L
x9L
x8L
x7L
x6L
x5L
x4L
x3L
x2L
x1L
x0L
x/L
x.L
x-L
x,L
x+L
x*L
x)L
x(L
x'L
0&L
0%L
0$L
0#L
0"L
0!L
0~K
0}K
0|K
0?M
0>M
x=M
x<M
x;M
x:M
x9M
x8M
x7M
x6M
x5M
x4M
x3M
x2M
x1M
x0M
x/M
x.M
x-M
x,M
x+M
x*M
x)M
x(M
x'M
x&M
x%M
x$M
x#M
x"M
x!M
x~L
x}L
x|L
x{L
xzL
xyL
xxL
xwL
xvL
xuL
xtL
xsL
xrL
xqL
0pL
0oL
0nL
0mL
0lL
0kL
0jL
0iL
0hL
0gL
0fL
0eL
0dL
0cL
0bL
0aL
0`L
0_L
0^L
0!N
0~M
0}M
0|M
0{M
0zM
0yM
0xM
0wM
xvM
xuM
xtM
xsM
xrM
xqM
xpM
xoM
xnM
xmM
xlM
xkM
xjM
xiM
xhM
xgM
xfM
xeM
xdM
xcM
xbM
xaM
x`M
x_M
x^M
x]M
x\M
x[M
xZM
xYM
xXM
xWM
xVM
xUM
xTM
xSM
xRM
xQM
xPM
xOM
xNM
xMM
xLM
xKM
xJM
xIM
xHM
xGM
xFM
xEM
xDM
xCM
xBM
xAM
x@M
0aN
0`N
0_N
0^N
0]N
0\N
0[N
0ZN
0YN
0XN
0WN
0VN
0UN
0TN
0SN
0RN
0QN
0PN
0ON
0NN
0MN
xLN
xKN
xJN
xIN
xHN
xGN
xFN
xEN
xDN
xCN
xBN
xAN
x@N
x?N
x>N
x=N
x<N
x;N
x:N
x9N
x8N
x7N
x6N
x5N
x4N
x3N
x2N
x1N
x0N
x/N
x.N
x-N
x,N
x+N
x*N
x)N
x(N
x'N
x&N
x%N
x$N
x#N
x"N
xCO
xBO
xAO
x@O
x?O
x>O
x=O
x<O
x;O
x:O
x9O
x8O
x7O
x6O
x5O
x4O
x3O
x2O
x1O
x0O
x/O
x.O
x-O
x,O
x+O
x*O
x)O
x(O
x'O
x&O
x%O
x$O
x#O
x"O
x!O
x~N
x}N
x|N
x{N
xzN
xyN
xxN
xwN
xvN
xuN
xtN
xsN
xrN
xqN
xpN
xoN
xnN
xmN
xlN
xkN
xjN
xiN
xhN
xgN
xfN
xeN
xdN
xcN
xbN
0%P
x$P
x#P
x"P
x!P
x~O
x}O
x|O
x{O
xzO
xyO
xxO
xwO
xvO
xuO
xtO
xsO
xrO
xqO
xpO
xoO
xnO
xmO
xlO
xkO
xjO
xiO
xhO
xgO
xfO
xeO
xdO
xcO
xbO
xaO
x`O
x_O
x^O
x]O
x\O
x[O
xZO
xYO
xXO
xWO
xVO
xUO
xTO
xSO
xRO
xQO
xPO
xOO
xNO
xMO
xLO
xKO
xJO
xIO
xHO
xGO
xFO
xEO
xDO
0eP
xdP
xcP
xbP
xaP
x`P
x_P
x^P
x]P
x\P
x[P
xZP
xYP
xXP
xWP
xVP
xUP
xTP
xSP
xRP
xQP
xPP
xOP
xNP
xMP
xLP
xKP
xJP
xIP
xHP
xGP
xFP
xEP
xDP
xCP
xBP
xAP
x@P
x?P
x>P
x=P
x<P
x;P
x:P
x9P
x8P
x7P
x6P
x5P
x4P
x3P
x2P
x1P
x0P
x/P
x.P
0-P
0,P
0+P
0*P
0)P
0(P
0'P
0&P
xGQ
xFQ
xEQ
xDQ
xCQ
xBQ
xAQ
x@Q
x?Q
x>Q
x=Q
x<Q
x;Q
x:Q
x9Q
x8Q
x7Q
x6Q
x5Q
x4Q
x3Q
x2Q
x1Q
x0Q
x/Q
x.Q
x-Q
x,Q
x+Q
x*Q
x)Q
x(Q
x'Q
x&Q
x%Q
x$Q
x#Q
x"Q
x!Q
x~P
x}P
x|P
x{P
xzP
xyP
xxP
xwP
xvP
xuP
xtP
xsP
xrP
xqP
xpP
xoP
0nP
0mP
0lP
0kP
0jP
0iP
0hP
0gP
0fP
x$W
x#W
x"W
x!W
x~V
x}V
x|V
x{V
xzV
xyV
xxV
xwV
xvV
xuV
xtV
xsV
xrV
xqV
xpV
xoV
xnV
xmV
xlV
xkV
xjV
xiV
xhV
xgV
xfV
xeV
xdV
xcV
xbV
xaV
x`V
x_V
x^V
x]V
x\V
x[V
xZV
xYV
xXV
xWV
xVV
xUV
xTV
xSV
xRV
xQV
xPV
xOV
xNV
xMV
xLV
0KV
0JV
0IV
0HV
0GV
0FV
0EV
0DV
0CV
0dW
0cW
0bW
0aW
0`W
0_W
0^W
0]W
0\W
x[W
xZW
xYW
xXW
xWW
xVW
xUW
xTW
xSW
xRW
xQW
xPW
xOW
xNW
xMW
xLW
xKW
xJW
xIW
xHW
xGW
xFW
xEW
xDW
xCW
xBW
xAW
x@W
x?W
x>W
x=W
x<W
x;W
x:W
x9W
x8W
x7W
x6W
x5W
x4W
x3W
x2W
x1W
x0W
x/W
x.W
x-W
x,W
x+W
x*W
x)W
x(W
x'W
x&W
x%W
xFX
xEX
xDX
xCX
xBX
xAX
x@X
x?X
x>X
x=X
x<X
x;X
x:X
x9X
x8X
x7X
x6X
x5X
x4X
x3X
x2X
x1X
x0X
x/X
x.X
x-X
x,X
x+X
x*X
x)X
x(X
x'X
x&X
x%X
x$X
x#X
x"X
x!X
x~W
x}W
x|W
x{W
xzW
xyW
xxW
xwW
xvW
xuW
xtW
xsW
xrW
xqW
xpW
xoW
xnW
xmW
xlW
xkW
xjW
xiW
xhW
xgW
xfW
xeW
xjY
xiY
xhY
xgY
xfY
xeY
xdY
xcY
xbY
xaY
x`Y
x_Y
x^Y
x]Y
x\Y
x[Y
xZY
xYY
xXY
xWY
xVY
xUY
xTY
xSY
xRY
xQY
xPY
xOY
xNY
xMY
xLY
xKY
xJY
xIY
xHY
xGY
xFY
xEY
xDY
xCY
xBY
xAY
x@Y
x?Y
x>Y
x=Y
x<Y
x;Y
x:Y
x9Y
x8Y
x7Y
x6Y
x5Y
x4Y
x3Y
x2Y
x1Y
x0Y
x/Y
x.Y
x-Y
x,Y
x+Y
x*Y
0)Y
0(Y
0'Y
0&Y
0%Y
0$Y
0#Y
0"Y
0!Y
0~X
0}X
0|X
0{X
0zX
0yX
0xX
0wX
0vX
0uX
0tX
0sX
0rX
0qX
0pX
0oX
0nX
0mX
0lX
0kX
0jX
0iX
0hX
0gX
0fX
0eX
0dX
0cX
0bX
0aX
0`X
0_X
0^X
0]X
0\X
0[X
0ZX
0YX
0XX
0WX
0VX
0UX
0TX
0SX
0RX
0QX
0PX
0OX
0NX
0MX
0LX
0KX
0JX
0IX
0HX
0u!
0t!
0s!
0r!
0q!
0p!
0o!
0n!
0m!
0l!
0k!
0j!
0i!
0h!
0g!
0f!
0e!
0d!
0c!
0b!
0a!
0`!
0_!
0^!
0]!
0\!
0[!
0Z!
0Y!
0X!
0W!
0V!
07"
06"
05"
04"
03"
02"
01"
00"
0/"
0."
0-"
0,"
0+"
0*"
0)"
0("
0'"
0&"
0%"
0$"
0#"
0""
0!"
0~!
0}!
0|!
0{!
0z!
0y!
0x!
0w!
0v!
1U!
0T!
0JQ
$end
#1800
1"
1T!
b0 N:
b100000000000000000000000000000000000 O:
b1010100000000000000000000000000000000000 P:
b0 Q:
b1010100000000000000000000000000000000000 R:
b0 S:
b1010100000000000000000000000000000000000 T:
b0 U:
b1010100000000000000000000000000000000000 V:
b0 W:
b11110101010101010101010101010000000000 X:
b0 Y:
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx "F
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx0 #F
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx $F
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx0 %F
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 yK
bx0 zK
b0 P!
b0 H!
b0 I!
0vM
0=M
0*I
0)I
08G
0kF
0jF
04F
0$D
0#D
0"D
0!D
0~C
0}C
0|C
0{C
0zC
0yC
0xC
0wC
0vC
0uC
0tC
0sC
0rC
0qC
0pC
0oC
0nC
0mC
0lC
0kC
0jC
0iC
0hC
0gC
0fC
0eC
0dC
0cC
0bC
0aC
0`C
0YC
0XC
0WC
0VC
0UC
0TC
0SC
0RC
0QC
0PC
1OC
0NC
1MC
0LC
1KC
0JC
1IC
0HC
1GC
0FC
1EC
0DC
1CC
0BC
1AC
0@C
1?C
0>C
1=C
0<C
1;C
0:C
19C
08C
17C
16C
15C
14C
00C
0/C
0.C
0-C
0,C
0+C
0*C
0)C
0(C
0'C
0&C
0%C
0$C
0#C
0"C
0!C
0~B
0}B
0|B
0{B
0zB
0yB
0xB
0wB
0vB
0uB
0tB
0sB
0rB
0qB
0pB
0oB
0nB
0mB
0lB
0kB
0eB
0dB
0cB
0bB
0aB
0`B
0_B
0^B
0]B
0\B
0[B
0ZB
0YB
0XB
0WB
0VB
0UB
0TB
0SB
0RB
0QB
0PB
0OB
0NB
0MB
0LB
0KB
0JB
0IB
0HB
0GB
0FB
0EB
0DB
0CB
1BB
0AB
1@B
0?B
1>B
00@
0/@
0.@
0-@
0,@
0+@
0*@
0)@
0(@
0'@
0&@
0%@
0$@
0#@
0"@
0!@
0~?
0}?
0|?
0{?
0z?
0y?
0x?
0w?
0v?
0u?
0t?
0s?
0r?
0q?
0p?
0o?
0n?
0m?
0l?
0k?
0b?
0a?
0`?
0_?
0^?
0]?
0\?
0[?
0Z?
0Y?
0X?
0W?
0V?
0U?
0T?
0S?
0R?
0Q?
0P?
0O?
0N?
0M?
0L?
0K?
0J?
0I?
0H?
0G?
0F?
0E?
0D?
0C?
0B?
0A?
0@?
1??
0>?
1=?
0<?
1;?
06?
05?
04?
03?
02?
01?
00?
0/?
0.?
0-?
0,?
0+?
0*?
0)?
0(?
0'?
0&?
0%?
0$?
0#?
0"?
0!?
0~>
0}>
0|>
0{>
0z>
0y>
0x>
0w>
0v>
0u>
0t>
0s>
0r>
0q>
0h>
0g>
0f>
0e>
0d>
0c>
0b>
0a>
0`>
0_>
0^>
0]>
0\>
0[>
0Z>
0Y>
0X>
0W>
0V>
0U>
0T>
0S>
0R>
0Q>
0P>
0O>
0N>
0M>
0L>
0K>
0J>
0I>
0H>
0G>
0F>
1E>
0D>
1C>
0B>
1A>
0D<
0C<
0B<
0A<
0@<
0?<
0><
0=<
0<<
0;<
0:<
09<
08<
07<
06<
05<
04<
03<
02<
01<
00<
0/<
0.<
0-<
0,<
0+<
0*<
0)<
0(<
0'<
0&<
0%<
0$<
0#<
0"<
0!<
0z;
0y;
0x;
0w;
0v;
0u;
0t;
0s;
0r;
0q;
0p;
0o;
0n;
0m;
0l;
0k;
0j;
0i;
0h;
0g;
0f;
0e;
0d;
0c;
0b;
0a;
0`;
0_;
0^;
0];
0\;
0[;
0Z;
0Y;
0X;
1W;
0V;
1U;
0T;
1S;
0P;
0O;
0N;
0M;
0L;
0K;
0J;
0I;
0H;
0G;
0F;
0E;
0D;
0C;
0B;
0A;
0@;
0?;
0>;
0=;
0<;
0;;
0:;
09;
08;
07;
06;
05;
04;
03;
02;
01;
00;
0/;
0.;
1-;
0&;
0%;
0$;
0#;
0";
0!;
0~:
0}:
0|:
0{:
0z:
0y:
0x:
0w:
0v:
0u:
0t:
0s:
0r:
0q:
0p:
0o:
0n:
0m:
0l:
0k:
0j:
0i:
0h:
0g:
0f:
0e:
0d:
0c:
0b:
0a:
0NR
0MR
0LR
0KR
0JR
0IR
0HR
0GR
0FR
0ER
0DR
0CR
0BR
0AR
0@R
0?R
0>R
0=R
0<R
0;R
0:R
09R
08R
07R
06R
05R
04R
03R
02R
01R
00R
0/R
0.R
0-R
0,R
0+R
1*R
0A=
0@=
0?=
0>=
0==
0<=
0;=
0:=
09=
08=
07=
06=
05=
04=
03=
02=
01=
00=
0/=
0.=
0-=
0,=
0+=
0*=
0)=
0(=
0'=
0&=
0%=
0$=
0#=
0"=
0!=
0~<
0}<
0|<
0{<
0wR
0vR
0uR
0tR
0sR
0rR
0qR
0pR
0oR
0nR
0mR
0lR
0kR
0jR
0iR
0hR
0gR
0fR
0eR
0dR
0cR
0bR
0aR
0`R
0_R
0^R
0]R
0\R
0[R
0ZR
0YR
0XR
0WR
0VR
0UR
1TR
0SR
1RR
0QR
1PR
0q=
0p=
0o=
0vS
0uS
0tS
0sS
0rS
0qS
0pS
0oS
0nS
0mS
0lS
0kS
0jS
0iS
0hS
0gS
0fS
0eS
0dS
0cS
0bS
0aS
0`S
0_S
0^S
0]S
0\S
0[S
0ZS
0YS
0XS
0WS
0VS
0US
0TS
1SS
0RS
1QS
0PS
1OS
09A
08A
07A
06A
05A
04A
03A
02A
01A
00A
0/A
0.A
0-A
0,A
0+A
0*A
0)A
0(A
0'A
0&A
0%A
0$A
0#A
0"A
0!A
0~@
0}@
0|@
0{@
0z@
0y@
0x@
0w@
0v@
0u@
0s@
0q@
0AT
0@T
0?T
0>T
0=T
0<T
0;T
0:T
09T
08T
07T
06T
05T
04T
03T
02T
01T
00T
0/T
0.T
0-T
0,T
0+T
0*T
0)T
0(T
0'T
0&T
0%T
0$T
0#T
0"T
0!T
0~S
0}S
1|S
0{S
1zS
0yS
1xS
0nA
0mA
0lA
0kA
0EU
0DU
0CU
0BU
0AU
0@U
0?U
0>U
0=U
0<U
0;U
0:U
09U
08U
07U
06U
05U
04U
03U
02U
01U
00U
0/U
0.U
0-U
0,U
0+U
0*U
0)U
0(U
0'U
0&U
0%U
0$U
0#U
1"U
0!U
1~T
0}T
1|T
0'E
0&E
0%E
0$E
0#E
0"E
0!E
0~D
0}D
0|D
0{D
0zD
0yD
0xD
0wD
0vD
0tD
0rD
0pD
0nD
0lD
0jD
0hD
0fD
0dD
0kU
0jU
0iU
0hU
0gU
0fU
0eU
0dU
0cU
0bU
1aU
0`U
1_U
0^U
1]U
0\U
1[U
0ZU
1YU
0XU
1WU
0VU
1UU
0TU
1SU
0RU
1QU
0PU
1OU
0NU
1MU
0LU
1KU
0JU
1IU
1HU
1GU
1FU
0VE
0UE
0TE
0oG
0TH
0SH
0[W
0XD
0WD
0VD
0UD
0TD
0SD
0RD
0QD
0PD
0OD
0ND
0MD
0LD
0KD
0JD
0ID
0GD
0ED
0CD
0AD
0?D
0=D
0;D
09D
07D
0?V
0>V
0=V
0<V
0;V
0:V
09V
08V
07V
06V
05V
04V
03V
02V
01V
00V
1/V
0.V
1-V
0,V
1+V
0*V
1)V
0(V
1'V
0&V
1%V
0$V
1#V
0"V
1!V
0~U
1}U
0|U
1{U
1zU
1yU
1xU
1wU
1vU
1uU
1tU
1sU
1rU
0uD
0sD
0qD
0oD
0mD
0kD
0iD
0gD
0eD
0cD
0bD
0aD
0`D
0_D
0^D
0g@
0f@
0e@
0d@
0c@
0b@
0a@
0`@
0_@
0^@
0]@
0\@
0[@
0Z@
0Y@
0X@
0W@
0V@
0U@
0T@
0S@
0R@
0Q@
0P@
0O@
0N@
0M@
0L@
0K@
0J@
0I@
0H@
0G@
0F@
0E@
0C@
0A@
0vT
0uT
0tT
0sT
0rT
0qT
0pT
0oT
0nT
0mT
0lT
0kT
0jT
0iT
0hT
0gT
0fT
0eT
0dT
0cT
0bT
0aT
0`T
0_T
0^T
0]T
0\T
0[T
0ZT
0YT
0XT
0WT
0VT
0UT
0TT
1ST
0RT
1QT
0PT
1OT
0NT
1MT
0LT
1KT
0JT
1IT
0t@
0r@
0p@
0s<
0r<
0q<
0p<
0o<
0n<
0m<
0l<
0k<
0j<
0i<
0h<
0g<
0f<
0e<
0d<
0c<
0b<
0a<
0`<
0_<
0^<
0]<
0\<
0[<
0Z<
0Y<
0X<
0W<
0V<
0U<
0T<
0S<
0R<
0Q<
0P<
0O<
0FS
0ES
0DS
0CS
0BS
0AS
0@S
0?S
0>S
0=S
0<S
0;S
0:S
09S
08S
07S
06S
05S
04S
03S
02S
01S
00S
0/S
0.S
0-S
0,S
0+S
0*S
0)S
0(S
0'S
0&S
0%S
0$S
0#S
1"S
1!S
0~R
1}R
0|R
1{R
0l=
0k=
0j=
0i=
0h=
0g=
0f=
0e=
0d=
0c=
0b=
0a=
0`=
0_=
0^=
0]=
0\=
0[=
0Z=
0Y=
0X=
0W=
0V=
0U=
0T=
0S=
0R=
0Q=
0P=
0O=
0N=
0M=
0L=
0K=
0J=
0I=
1H=
1G=
0F=
1E=
0D=
1C=
08>
07>
06>
05>
04>
03>
02>
01>
00>
0/>
0.>
0->
0,>
0+>
0*>
0)>
0(>
0'>
0&>
0%>
0$>
0#>
0">
0!>
0~=
0}=
0|=
0{=
0z=
0y=
0x=
0w=
0v=
0u=
0t=
0s=
0r=
0D@
0B@
0@@
0hA
0gA
0fA
0eA
0dA
0cA
0bA
0aA
0`A
0_A
0^A
0]A
0\A
0[A
0ZA
0YA
0XA
0WA
0VA
0UA
0TA
0SA
0RA
0QA
0PA
0OA
0NA
0MA
0LA
0KA
0JA
0IA
0HA
0GA
0FA
1EA
1CA
1AA
1?A
0>A
1=A
0<A
1;A
08B
07B
06B
05B
04B
03B
02B
01B
00B
0/B
0.B
0-B
0,B
0+B
0*B
0)B
0(B
0'B
0&B
0%B
0$B
0#B
0"B
0!B
0~A
0}A
0|A
0{A
0zA
0yA
0xA
0wA
0vA
0uA
0tA
0sA
0rA
0qA
0pA
0oA
0HD
0FD
0DD
0BD
0@D
0>D
0<D
0:D
08D
06D
05D
04D
03D
02D
01D
0SE
0RE
0QE
0PE
0OE
0NE
0ME
0LE
0KE
0JE
0IE
0HE
0GE
0FE
0EE
0DE
1CE
1AE
1?E
1=E
1;E
19E
17E
15E
13E
11E
1*E
1)E
1(E
0~E
0}E
0|E
0{E
0zE
0yE
0xE
0wE
0vE
0uE
0tE
0sE
0rE
0qE
0pE
0oE
0nE
0mE
0lE
0kE
0jE
0iE
0hE
0gE
0fE
0eE
0dE
0cE
0bE
0aE
0`E
0_E
0^E
0]E
0BE
0@E
0>E
0<E
0:E
08E
06E
04E
02E
10E
1/E
1.E
1-E
1,E
1+E
0\E
0[E
0ZE
0YE
0XE
0WE
0DA
0BA
0@A
#3600
0"
0T!
#5400
1"
1T!
b101011000000000000000000000000000000000000 "F
b0 #F
b1010101010100000000000000000000000000000000000 $F
b0 %F
b11111111110101010101010101010000000000000000 &F
b0 'F
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx xK
b0xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00 yK
b0 Q!
b0 J!
b0 K!
0iY
0hY
0gY
0fY
0eY
0dY
0cY
0bY
0aY
0`Y
0_Y
0^Y
0]Y
0\Y
0[Y
0ZY
0YY
0XY
0WY
0VY
0UY
0TY
0SY
0RY
0QY
0PY
0OY
0NY
0MY
0LY
0KY
0JY
0IY
0HY
0GY
0FY
0EY
0DY
0CY
0BY
0AY
0@Y
0?Y
0>Y
0=Y
0<Y
0;Y
0:Y
09Y
08Y
07Y
06Y
05Y
04Y
03Y
02Y
01Y
00Y
0/Y
0.Y
0-Y
0,Y
0+Y
0*Y
0rL
0qL
0'L
0ZJ
0YJ
0XJ
0WJ
0VJ
0UJ
0TJ
0SJ
0RJ
0QJ
0PJ
0OJ
0NJ
0MJ
0LJ
0KJ
0JJ
0IJ
0HJ
0GJ
0FJ
0EJ
0DJ
0CJ
0BJ
0AJ
0@J
0?J
0>J
0=J
0<J
0;J
0:J
09J
08J
07J
06J
05J
04J
03J
02J
01J
0%J
0$J
0#J
0"J
0!J
0~I
0}I
0|I
0{I
0zI
0yI
0xI
0wI
0vI
0uI
0tI
1sI
0rI
1qI
0pI
1oI
0nI
1mI
0lI
1kI
0jI
1iI
0hI
1gI
0fI
1eI
0dI
1cI
0bI
1aI
1`I
1_I
1^I
1]I
1\I
1[I
1ZI
1YI
1XI
0VI
0UI
0TI
0SI
0RI
0QI
0PI
0OI
0NI
0MI
0LI
0KI
0JI
0II
0HI
0GI
0FI
0EI
0DI
0CI
0BI
0AI
0@I
0?I
0>I
0=I
0<I
0;I
0:I
09I
08I
07I
06I
05I
04I
03I
02I
01I
00I
0/I
0.I
0-I
0,I
0+I
0fG
0eG
0dG
0cG
0bG
0aG
0`G
0_G
0^G
0]G
0\G
0[G
0ZG
0YG
0XG
0WG
0VG
0UG
0TG
0SG
0RG
0QG
0PG
0OG
0NG
0MG
0LG
0KG
0JG
0IG
0HG
0GG
0FG
0EG
0DG
1CG
0BG
1AG
0@G
1?G
0>G
1=G
0<G
1;G
0:G
19G
05G
04G
03G
02G
01G
00G
0/G
0.G
0-G
0,G
0+G
0*G
0)G
0(G
0'G
0&G
0%G
0$G
0#G
0"G
0!G
0~F
0}F
0|F
0{F
0zF
0yF
0xF
0wF
0vF
0uF
0tF
0sF
0rF
0qF
0pF
0oF
0nF
0mF
0lF
0^F
0]F
0\F
0[F
0ZF
0YF
0XF
0WF
0VF
0UF
0TF
0SF
0RF
0QF
0PF
0OF
0NF
0MF
0LF
0KF
0JF
0IF
0HF
0GF
0FF
0EF
0DF
0CF
0BF
0AF
0@F
0?F
0>F
0=F
0<F
0;F
1:F
19F
08F
17F
06F
15F
0GH
0FH
0EH
0DH
0CH
0BH
0AH
0@H
0?H
0>H
0=H
0<H
0;H
0:H
09H
08H
07H
06H
05H
04H
03H
02H
01H
00H
0/H
0.H
0-H
0,H
0+H
0*H
0)H
0(H
0'H
0&H
0%H
0$H
1#H
1"H
0!H
1~G
0}G
1|G
0{G
1zG
0yG
1xG
0wG
1vG
0uG
1tG
0sG
1rG
0qG
1pG
0|H
0{H
0zH
0yH
0xH
0wH
0vH
0uH
0tH
0sH
0rH
0qH
0pH
0oH
0nH
0mH
0lH
0kH
0jH
0iH
0hH
0gH
0fH
0eH
0dH
0cH
0bH
0aH
0`H
0_H
0^H
0]H
0\H
0[H
0ZH
0YH
0XH
0WH
0VH
0UH
0?K
0>K
0=K
0<K
0;K
0:K
09K
08K
07K
06K
05K
04K
03K
02K
01K
00K
0/K
0.K
0-K
0,K
0+K
0*K
0)K
0(K
0'K
0&K
1%K
0$K
1#K
0"K
1!K
0~J
1}J
0|J
1{J
0zJ
1yJ
0xJ
1wJ
0vJ
1uJ
0tJ
1sJ
0rJ
1qJ
1pJ
1oJ
1nJ
1mJ
1lJ
1kJ
1jJ
1iJ
1hJ
0lK
0kK
0jK
0iK
0hK
0gK
0fK
0eK
0dK
0cK
0bK
0aK
0`K
0_K
0^K
0]K
0\K
0[K
0ZK
0YK
0XK
0WK
0VK
0UK
0TK
0SK
0RK
0QK
0PK
0OK
0NK
0MK
0LK
0KK
0JK
0IK
0HK
0GK
0FK
0EK
0DK
0CK
0BK
0AK
0LV
0oP
0.P
#7200
0"
0T!
#9000
1"
1T!
b101010101010101011000000000000000000000000000000000000 xK
b0 yK
b1111111111010101010101010101000000000000000000000000000 zK
b0 {K
b0 R!
b0 L!
b0 M!
0LN
0KN
0JN
0IN
0HN
0GN
0FN
0EN
0DN
0CN
0BN
0AN
0@N
0?N
0>N
0=N
0<N
0;N
0:N
09N
08N
07N
06N
05N
04N
03N
02N
01N
00N
0/N
0.N
0-N
0,N
0+N
0*N
0)N
0(N
0'N
0&N
0%N
0$N
0#N
0"N
0uM
0tM
0sM
0rM
0qM
0pM
0oM
0nM
0mM
0lM
0kM
0jM
0iM
0hM
0gM
0fM
0eM
0dM
0cM
0bM
0aM
0`M
0_M
0^M
0]M
0\M
1[M
0ZM
1YM
0XM
1WM
0VM
1UM
0TM
1SM
0RM
1QM
0PM
1OM
0NM
1MM
0LM
1KM
0JM
1IM
1HM
1GM
1FM
1EM
1DM
1CM
1BM
1AM
1@M
0<M
0;M
0:M
09M
08M
07M
06M
05M
04M
03M
02M
01M
00M
0/M
0.M
0-M
0,M
0+M
0*M
0)M
0(M
0'M
0&M
0%M
0$M
0#M
0"M
0!M
0~L
0}L
0|L
0{L
0zL
0yL
0xL
0wL
0vL
0uL
0tL
0sL
0]L
0\L
0[L
0ZL
0YL
0XL
0WL
0VL
0UL
0TL
0SL
0RL
0QL
0PL
0OL
0NL
0ML
0LL
0KL
0JL
0IL
0HL
0GL
0FL
0EL
0DL
0CL
0BL
0AL
0@L
0?L
0>L
0=L
0<L
0;L
0:L
19L
18L
07L
16L
05L
14L
03L
12L
01L
10L
0/L
1.L
0-L
1,L
0+L
1*L
0)L
1(L
0$W
0#W
0"W
0!W
0~V
0}V
0|V
0{V
0zV
0yV
0xV
0wV
0vV
0uV
0tV
0sV
0rV
0qV
0pV
0oV
0nV
0mV
0lV
0kV
0jV
0iV
0hV
0gV
0fV
0eV
0dV
0cV
0bV
0aV
0`V
0_V
1^V
1]V
0\V
1[V
0ZV
1YV
0XV
1WV
0VV
1UV
0TV
1SV
0RV
1QV
0PV
1OV
0NV
1MV
0GQ
0FQ
0EQ
0DQ
0CQ
0BQ
0AQ
0@Q
0?Q
0>Q
0=Q
0<Q
0;Q
0:Q
09Q
08Q
07Q
06Q
05Q
04Q
03Q
02Q
01Q
00Q
0/Q
0.Q
0-Q
0,Q
0+Q
0*Q
0)Q
0(Q
0'Q
0&Q
0%Q
0$Q
0ZW
0YW
0XW
0WW
0VW
0UW
0TW
0SW
0RW
0QW
0PW
0OW
0NW
0MW
0LW
0KW
0JW
0IW
0HW
0GW
0FW
0EW
0DW
0CW
0BW
0AW
1@W
0?W
1>W
0=W
1<W
0;W
1:W
09W
18W
07W
16W
05W
14W
03W
12W
01W
10W
0/W
1.W
1-W
1,W
1+W
1*W
1)W
1(W
1'W
1&W
1%W
0LO
0KO
0JO
0IO
0HO
0GO
0FO
0EO
0DO
0dP
0cP
0bP
0aP
0`P
0_P
0^P
0]P
0\P
0[P
0ZP
0YP
0XP
0WP
0VP
0UP
0TP
0SP
0RP
0QP
0PP
0OP
0NP
0MP
0LP
0KP
0JP
0IP
0HP
0GP
0FP
0EP
0DP
0CP
0BP
0AP
0FX
0EX
0DX
0CX
0BX
0AX
0@X
0?X
0>X
0=X
0<X
0;X
0:X
09X
08X
07X
06X
05X
04X
03X
02X
01X
00X
0/X
0.X
0-X
0,X
0+X
0*X
0)X
0(X
0'X
0&X
0%X
0$X
0#X
0"X
1!X
1~W
1}W
1|W
1{W
1zW
1yW
1xW
1wW
1vW
1uW
1tW
1sW
1rW
1qW
1pW
1oW
1nW
1mW
1lW
1kW
1jW
1iW
1hW
1gW
1fW
1eW
1#Q
0"Q
0!Q
0~P
0}P
0|P
0{P
0zP
0yP
0xP
0wP
0vP
0uP
0tP
0sP
0rP
0qP
0pP
1@P
0?P
0>P
0=P
0<P
0;P
0:P
09P
08P
07P
06P
05P
04P
03P
02P
01P
00P
0/P
0CO
0BO
0AO
0@O
0?O
0>O
0=O
0<O
0;O
0:O
09O
08O
07O
06O
05O
04O
03O
02O
01O
00O
0/O
0.O
0-O
0,O
0+O
0*O
0)O
0(O
0'O
0&O
0%O
0$O
0#O
0"O
0!O
0~N
0}N
1jN
1iN
1hN
1gN
1fN
1eN
1dN
1cN
1bN
0$P
0#P
0"P
0!P
0~O
0}O
0|O
0{O
0zO
0yO
0xO
0wO
0vO
0uO
0tO
0sO
0rO
0qO
0pO
0oO
0nO
0mO
0lO
0kO
0jO
0iO
0hO
0gO
0fO
0eO
0dO
0cO
0bO
0aO
0`O
0_O
0|N
1{N
1zN
1yN
1xN
1wN
1vN
1uN
1tN
1sN
1rN
1qN
1pN
1oN
1nN
1mN
1lN
1kN
1^O
0]O
0\O
0[O
0ZO
0YO
0XO
0WO
0VO
0UO
0TO
0SO
0RO
0QO
0PO
0OO
0NO
0MO
#10800
0"
0T!
#12600
1"
1T!
b1111111111111111111111111100000000000000000000000000000000000000 HQ
b10000000000000000000000000000000000000 IQ
b0 S!
b0 N!
b0 O!
0c
0b
0a
0`
0_
0^
0]
0\
0[
0Z
0Y
0X
0W
0V
0U
0T
0S
0R
0Q
0P
0O
0N
0M
0L
0K
0J
0I
0H
0G
0F
0E
0D
0C
0B
0A
0@
0?
0>
0=
0<
0;
0:
09
08
07
06
05
04
03
02
01
00
0/
0.
0-
0,
0+
0*
0)
0(
0'
0&
0%
0$
1jY
#14400
0"
0T!
#16200
1"
1T!
#18000
0"
0T!
#19800
1"
1T!
#21600
0"
0T!
#23400
1"
1T!
#25200
0"
0T!
#27000
1"
1T!
#28800
0"
0T!
#30600
1"
1T!
#32400
0"
0T!
#34200
1"
1T!
#36000
0"
0T!
#37800
1"
1T!
#39600
b10010000101010011010100100100 d
b11000000100010010101111010000001 e
0"
1)Y
1"Y
1~X
1}X
1|X
1{X
1yX
1wX
1tX
1pX
1iX
1hX
1u!
1n!
1l!
1k!
1j!
1i!
1g!
1e!
1b!
1^!
1W!
1V!
1eX
1bX
1_X
1]X
1[X
1ZX
1WX
1UX
1SX
1NX
1KX
1E!
1B!
1?!
1>!
1=!
1<!
1;!
1:!
19!
18!
16!
15!
13!
12!
11!
1.!
1-!
1+!
1)!
1'!
1%!
1$!
1#!
1"!
1~
1|
1{
1x
1w
1s
1n
1m
1l
1j
1i
1h
1g
1f
0T!
1r(
1k(
1i(
1h(
1g(
1f(
1d(
1b(
1_(
1[(
1T(
1S(
15"
12"
1/"
1-"
1+"
1*"
1'"
1%"
1#"
1|!
1y!
b1 pQ
b1 ^Q
b1 RQ
0PQ
0VQ
0YQ
0\Q
0bQ
0eQ
0hQ
0kQ
0tQ
0wQ
b111000000100010010101111010000001 NQ
b1111110111011010100001011111101 QQ
b111000000100010010101111010000001 TQ
b111000000100010010101111010000001 WQ
b111000000100010010101111010000001 ZQ
b111111011101101010000101111110 ]Q
b111000000100010010101111010000001 `Q
b111000000100010010101111010000001 cQ
b111000000100010010101111010000001 fQ
b111000000100010010101111010000001 iQ
b1111110111011010100001011111101 oQ
b111000000100010010101111010000001 rQ
b111000000100010010101111010000001 uQ
0$)
0")
0!)
0~(
0|(
0{(
0z(
0y(
0v(
0u(
1P'
1I'
1G'
1F'
1E'
1D'
1B'
1@'
1='
19'
12'
11'
10'
1/'
1('
1&'
1%'
1$'
1#'
1!'
1}&
1z&
1v&
1o&
1n&
1m&
1l&
1j&
1i&
1h&
1g&
1f&
1e&
1c&
1^&
1\&
1Z&
1Y&
1W&
1V&
1U&
1S&
1R&
1Q&
1P&
1O&
1N&
1*&
1#&
1!&
1~%
1}%
1|%
1z%
1x%
1u%
1q%
1j%
1i%
1h%
1g%
1`%
1^%
1]%
1\%
1[%
1Y%
1W%
1T%
1P%
1I%
1H%
1G%
1F%
1?%
1=%
1<%
1;%
1:%
18%
16%
13%
1/%
1(%
1'%
1&%
1%%
1|$
1z$
1y$
1x$
1w$
1u$
1s$
1p$
1l$
1e$
1d$
1c$
1a$
1`$
1_$
1^$
1]$
1\$
1Z$
1U$
1S$
1Q$
1P$
1N$
1M$
1L$
1J$
1I$
1H$
1G$
1F$
1E$
1A$
1:$
18$
17$
16$
15$
13$
11$
1.$
1*$
1#$
1"$
1!$
1~#
1w#
1u#
1t#
1s#
1r#
1p#
1n#
1k#
1g#
1`#
1_#
1^#
1]#
1V#
1T#
1S#
1R#
1Q#
1O#
1M#
1J#
1F#
1?#
1>#
1=#
1<#
1:#
19#
18#
17#
16#
15#
13#
1.#
1,#
1*#
1)#
1'#
1&#
1%#
1##
1"#
1!#
1~"
1}"
1|"
1y"
1r"
1p"
1o"
1n"
1m"
1k"
1i"
1f"
1b"
1["
1Z"
1Y"
18(
1@(
1L(
1-,
1+,
1*,
1),
1(,
1',
1&,
1$,
1}+
1{+
1y+
1x+
1v+
1u+
1t+
1r+
1q+
1p+
1o+
1n+
1m+
1P/
1O/
1N/
1M/
1L/
1K/
1I/
1D/
1B/
1@/
1?/
1=/
1</
1;/
19/
18/
17/
16/
15/
14/
1M5
1K5
1J5
1I5
1H5
1G5
1F5
1D5
1?5
1=5
1;5
1:5
185
175
165
145
135
125
115
105
1/5
1#8
1z7
1x7
1w7
1v7
1u7
1s7
1q7
1n7
1j7
1c7
1b7
1a7
0`7
1u5
1s5
1l5
1j5
1i5
1h5
1g5
1e5
1c5
1`5
1\5
1U5
1T5
1S5
0R5
1u2
1n2
1l2
1k2
1j2
1i2
1g2
1e2
1b2
1^2
1W2
1V2
1U2
0T2
1O2
1H2
1F2
1E2
1D2
1C2
1A2
1?2
1<2
182
112
102
1/2
0.2
1)2
1"2
1~1
1}1
1|1
1{1
1y1
1w1
1t1
1p1
1i1
1h1
1g1
0f1
1y/
1w/
1p/
1n/
1m/
1l/
1k/
1i/
1g/
1d/
1`/
1Y/
1X/
1W/
0V/
1+/
1$/
1"/
1!/
1~.
1}.
1{.
1y.
1v.
1r.
1k.
1j.
1i.
0h.
1y,
1r,
1p,
1o,
1n,
1m,
1k,
1i,
1f,
1b,
1[,
1Z,
1Y,
0X,
1U,
1S,
1L,
1J,
1I,
1H,
1G,
1E,
1C,
1@,
1<,
15,
14,
13,
02,
11*
1**
1(*
1'*
1&*
1%*
1#*
1!*
1|)
1x)
1q)
1p)
1o)
0n)
1?+
18+
16+
15+
14+
13+
11+
1/+
1,+
1(+
1!+
1~*
1}*
1|*
0B+
154
134
114
1.4
1+4
1*4
1'4
1&4
1%4
1"4
1!4
1~3
1z3
1x3
1u3
1t3
1o3
0n3
1T4
1R4
1Q4
1P4
1O4
1M4
1K4
1F4
1=4
1;4
1%:
1|9
1z9
0y9
1x9
0w9
0u9
0s9
1p9
1l9
0e9
1d9
0c9
0b9
1A:
1?:
1=:
1;:
1-:
1+:
1.7
1-7
1,7
1+7
1*7
1&7
1%7
1$7
1|6
1y6
1x6
1u6
1t6
1s6
1r6
1q6
1o6
0n6
1m6
0l6
1Y7
1W7
1P7
1K7
1I7
1G7
1D7
1@7
187
171
151
141
121
111
1/1
1.1
1+1
1*1
1&1
1%1
1!1
1~0
1}0
1{0
1y0
1x0
1u0
0t0
1s0
0r0
1q0
0p0
1[1
1X1
1U1
1T1
1Q1
1P1
1O1
1L1
1K1
1H1
1D1
1A1
1@1
1<1
16.
14.
13.
12.
1-.
1+.
1*.
1).
1'.
1&.
1%.
1#.
1}-
1{-
1z-
1y-
1w-
0v-
1s-
0r-
1a.
1_.
1].
1X.
1V.
1T.
1S.
1Q.
1O.
1L.
1J.
1H.
1F.
1@.
1?.
#41400
1"
1T!
b111100000010001001010111101000000100 N:
b0 O:
b110010111010001011101110100001110100000 P:
b1100000101010100101011010100001010100 Q:
b101010011010111000110001100110110110100 R:
b10001100100010011001110011001001000000 S:
b110101100101000111001110011001001010100 T:
b1010000000010000101011110100000000000 U:
b101111111001100100000111000111110000000 V:
b10000000100010010101000010000001010000 W:
b11001001010111011100000010111000000100 X:
b10100000000000001010101000000000000 Y:
b1111101110000100011001101011110101010110011101101111111100100100 P!
b10010000101010011010100100100 H!
b11000000100010010101111010000001 I!
1xC
1vC
1tC
1rC
1dC
1bC
1WC
1PC
1NC
0MC
1LC
0KC
0IC
0GC
1DC
1@C
09C
18C
07C
06C
1.C
1,C
1%C
1~B
1|B
1zB
1wB
1sB
1kB
1^B
1]B
1\B
1[B
1ZB
1VB
1UB
1TB
1NB
1KB
1JB
1GB
1FB
1EB
1DB
1CB
1AB
0@B
1?B
0>B
1'@
1%@
1$@
1#@
1"@
1~?
1|?
1w?
1n?
1l?
1`?
1^?
1\?
1Y?
1V?
1U?
1R?
1Q?
1P?
1M?
1L?
1K?
1G?
1E?
1B?
1A?
1<?
0;?
12?
1/?
1,?
1+?
1(?
1'?
1&?
1#?
1"?
1}>
1y>
1v>
1u>
1q>
1f>
1d>
1c>
1a>
1`>
1^>
1]>
1Z>
1Y>
1U>
1T>
1P>
1O>
1N>
1L>
1J>
1I>
1F>
0E>
1D>
0C>
1B>
0A>
1D<
1B<
1@<
1;<
19<
17<
16<
14<
12<
1/<
1-<
1+<
1)<
1#<
1"<
1u;
1s;
1r;
1q;
1l;
1j;
1i;
1h;
1f;
1e;
1d;
1b;
1^;
1\;
1[;
1Z;
1X;
0W;
1T;
0S;
0-;
1$;
1{:
1y:
1x:
1w:
1v:
1t:
1r:
1o:
1k:
1d:
1c:
1b:
1a:
1LR
1ER
1CR
1BR
1AR
1@R
1>R
1<R
19R
15R
1.R
1-R
1,R
1+R
0*R
1?=
18=
16=
15=
14=
13=
11=
1/=
1,=
1(=
1!=
1~<
1}<
1|<
1{<
1tR
1oR
1nR
1kR
1eR
1dR
1cR
1aR
1]R
1XR
1WR
1UR
0TR
1SR
0RR
1QR
0PR
14>
12>
10>
1+>
1)>
1'>
1&>
1$>
1">
1}=
1{=
1y=
1w=
1q=
1tS
1rS
1qS
1nS
1kS
1iS
1gS
1eS
1dS
1bS
1`S
1_S
1^S
1]S
1ZS
1WS
1US
0SS
1RS
0QS
0OS
17A
15A
14A
12A
11A
1/A
1.A
1+A
1*A
1&A
1%A
1!A
1~@
1}@
1{@
1y@
1x@
1u@
1t@
1s@
1q@
1p@
1?T
1=T
1;T
18T
14T
13T
12T
1/T
1.T
1+T
1*T
1'T
1&T
1$T
1!T
1~S
0|S
0zS
1yS
0xS
1'B
1%B
1$B
1#B
1"B
1~A
1|A
1wA
1@U
1=U
1<U
1;U
1:U
17U
16U
15U
14U
12U
10U
1*U
1&U
1%U
1$U
1#U
1!U
0~T
0|T
1~D
1}D
1|D
1{D
1zD
1vD
1uD
1tD
1nD
1kD
1jD
1gD
1fD
1eD
1dD
1cD
1aD
1_D
1^D
1iU
1bU
1`U
0_U
0]U
1\U
0[U
1ZU
0YU
1XU
1VU
1RU
0KU
0IU
1lE
1jE
1hE
1fE
1QD
1PD
1OD
1ND
1MD
1ID
1HD
1GD
1AD
1>D
1=D
1:D
19D
18D
17D
16D
14D
12D
11D
1:V
16V
15V
14V
11V
0/V
0-V
1,V
0+V
0)V
1(V
0'V
1&V
0}U
1|U
0{U
0yU
0xU
0wU
0vU
0uU
0|D
0{D
0zD
1rD
0dD
0^D
1e@
1c@
1b@
1`@
1_@
1]@
1\@
1Y@
1X@
1T@
1S@
1O@
1N@
1M@
1K@
1I@
1H@
1E@
1D@
1C@
1A@
1@@
1tT
1rT
1qT
1lT
1kT
1jT
1iT
1eT
1dT
1cT
1aT
1`T
1_T
1YT
1WT
1VT
1RT
0QT
1PT
0MT
0KT
1JT
0IT
07A
05A
04A
0.A
1'A
0%A
1#A
1"A
0~@
0x@
1v@
0t@
0s@
0p@
1q<
1j<
1h<
1g<
1f<
1e<
1c<
1a<
1^<
1Z<
1S<
1R<
1Q<
1P<
1O<
1DS
1AS
1=S
1<S
1:S
19S
16S
14S
12S
10S
1.S
1-S
1*S
1&S
1#S
0!S
1~R
0}R
1|R
0{R
0?=
05=
04=
03=
0,=
0(=
0|<
0{<
0q<
0g<
0f<
0e<
0^<
0Z<
0P<
0O<
1j=
1i=
1g=
1c=
1^=
1]=
1\=
1[=
1Z=
1Y=
1X=
1T=
1S=
1R=
1P=
1L=
1K=
1J=
0H=
1F=
0E=
1D=
0C=
04>
00>
1/>
1->
1,>
0)>
0'>
1#>
0{=
0w=
1t=
1s=
0q=
1p=
0e@
0c@
0b@
0\@
1U@
0S@
1Q@
1P@
0N@
0H@
1F@
0D@
0C@
0@@
1fA
1eA
1dA
1bA
1`A
1_A
1^A
1[A
1YA
1XA
1WA
1VA
1UA
1TA
1RA
1QA
1OA
1NA
1MA
0EA
1BA
0AA
1@A
0?A
0=A
1<A
0;A
14B
1.B
1-B
0'B
0#B
0"B
1zA
1xA
1tA
1sA
1pA
1nA
1lA
0OD
0ND
0MD
1ED
07D
01D
1NE
1KE
1GE
1EE
1BE
1@E
0?E
0=E
1<E
1:E
18E
07E
14E
00E
0/E
0-E
1vE
1uE
1tE
0lE
0hE
0fE
1cE
1^E
1\E
1XE
1IE
1HE
0GE
1?E
01E
0+E
0uE
0tE
0eA
1cA
0bA
1\A
0UA
1SA
0QA
1PA
0NA
1HA
1FA
1DA
0CA
0@A
04B
0-B
1&B
0$B
1"B
0wA
0sA
0i=
1_=
0^=
0]=
1V=
0R=
1H=
0G=
0,>
0#>
0s=
#43200
b10000100100001001101011000001001 d
b10110001111100000101011001100011 e
0"
1(Y
1$Y
1#Y
0"Y
0|X
0wX
0tX
1sX
1rX
1qX
1oX
1kX
1jX
0iX
1t!
1p!
1o!
0n!
0j!
0e!
0b!
1a!
1`!
1_!
1]!
1Y!
1X!
0W!
1gX
0eX
1dX
0bX
0_X
1^X
0ZX
1YX
1XX
0WX
0SX
1PX
0NX
1MX
0KX
1HX
1G!
1F!
0E!
1D!
1C!
1A!
0=!
0;!
0:!
17!
06!
01!
10!
0.!
0-!
0+!
1(!
0'!
0%!
0$!
0"!
1!!
0|
1y
0x
0w
1u
1t
1p
0l
1k
0j
0i
0g
0f
0T!
1q(
1m(
1l(
0k(
0g(
0b(
0_(
1^(
1](
1\(
1Z(
1V(
1U(
0T(
17"
05"
14"
02"
0/"
1."
0*"
1)"
1("
0'"
0#"
1~!
0|!
1{!
0y!
1v!
b1 yQ
1wQ
b1 mQ
0qQ
b0 pQ
1kQ
0_Q
b0 ^Q
1bQ
b1 aQ
1YQ
b1 XQ
1VQ
0SQ
b0 RQ
1PQ
b1 OQ
0MQ
b110110001111100000101011001100011 KQ
b10011100000111110101001100111001 NQ
b110110001111100000101011001100011 QQ
b0 TQ
b10011100000111110101001100111001 WQ
b101100011111000001010110011000110 ZQ
b110110001111100000101011001100011 ]Q
b1001110000011111010100110011100 `Q
b110110001111100000101011001100011 cQ
b110110001111100000101011001100011 fQ
b0 iQ
b10011100000111110101001100111001 lQ
b110110001111100000101011001100011 oQ
b110110001111100000101011001100011 rQ
b0 uQ
b10011100000111110101001100111001 xQ
1u(
0w(
1y(
0}(
1|(
1!)
1")
0#)
1$)
0%)
1q'
1n'
1m'
1l'
1i'
1h'
1e'
1c'
1a'
1`'
1_'
1^'
1]'
1W'
1V'
1U'
1R'
0P'
0I'
0G'
0F'
0E'
0D'
0B'
0@'
0='
09'
02'
01'
00'
1.'
1*'
1)'
0('
0$'
0}&
0z&
1y&
1x&
1w&
1u&
1q&
1p&
0o&
1k&
0j&
0i&
0h&
0e&
1b&
1`&
0\&
0Z&
0Y&
1X&
1T&
0S&
0R&
0Q&
0N&
1M&
1L&
1K&
1H&
1G&
1F&
1C&
1B&
1?&
1=&
1;&
1:&
19&
18&
17&
11&
10&
1/&
1,&
0*&
0#&
0!&
0~%
0}%
0|%
0z%
0x%
0u%
0q%
0j%
0i%
0h%
1f%
1b%
1a%
0`%
0\%
0W%
0T%
1S%
1R%
1Q%
1O%
1K%
1J%
0I%
1E%
1A%
1@%
0?%
0;%
06%
03%
12%
11%
10%
1.%
1*%
1)%
0(%
0%%
1#%
1"%
1!%
1{$
0z$
0y$
0w$
1v$
0u$
1t$
1r$
1q$
0l$
1j$
1i$
1h$
0d$
0c$
1b$
0`$
0_$
0^$
0Z$
1Y$
1X$
1V$
0U$
1T$
0S$
0Q$
0P$
1K$
0I$
0H$
0G$
1C$
1B$
0A$
1@$
1?$
1;$
08$
05$
14$
03$
12$
01$
0.$
1,$
1+$
1)$
1($
1$$
0"$
1{#
1z#
1y#
0w#
1v#
0t#
0s#
1m#
1l#
1j#
0g#
1d#
1c#
1b#
0`#
0^#
0]#
0V#
0T#
0S#
0R#
0Q#
0O#
0M#
0J#
0F#
0?#
0>#
0=#
1;#
0:#
09#
08#
05#
12#
10#
0,#
0*#
0)#
1(#
1$#
0##
0"#
0!#
0|"
1{"
1z"
1v"
1u"
1t"
0r"
1q"
0o"
0n"
1h"
1g"
1e"
0b"
1_"
1^"
1]"
0["
0Y"
1X"
1W"
1S"
1R"
1O"
1N"
1L"
1J"
1D"
1C"
1B"
1A"
1@"
1<"
1;"
19"
18"
16(
08(
1<(
1B(
0@(
0L(
1J(
1R(
1m8
1-/
0+/
1*/
1)/
1%/
0"/
0}.
1|.
0{.
1z.
0y.
0v.
1t.
1s.
1q.
1p.
1l.
0j.
1+2
1(2
1$2
1#2
0"2
0|1
0w1
0t1
1s1
1r1
1q1
1o1
1k1
1j1
0i1
1N2
1J2
1I2
0H2
0D2
0?2
0<2
1;2
1:2
192
172
132
122
012
1'5
1$5
1#5
1"5
1}4
1|4
1y4
1w4
1u4
1t4
1s4
1r4
1q4
1k4
1j4
1i4
1f4
0u5
1r5
1n5
1m5
0l5
0h5
0c5
0`5
1_5
1^5
1]5
1[5
1W5
1V5
0U5
1G8
1D8
1C8
1B8
1?8
1>8
1;8
198
178
168
158
148
138
1-8
1,8
1+8
1(8
1m)
1l)
1h)
1g)
1d)
1c)
1a)
1_)
1Y)
1X)
1W)
1V)
1U)
1Q)
1P)
1N)
1M)
1L)
1K)
0J)
1.*
1-*
1,*
0**
1)*
0'*
0&*
1~)
1})
1{)
0x)
1u)
1t)
1s)
0q)
0o)
1n)
1/,
1,,
0+,
0*,
0),
0&,
1#,
1!,
0{+
0y+
0x+
1w+
1s+
0r+
0q+
0p+
0m+
1l+
1k+
0j+
0U,
0S,
0L,
0J,
0I,
0H,
0G,
0E,
0C,
0@,
0<,
05,
04,
03,
12,
1v,
1u,
1t,
0r,
1q,
0o,
0n,
1h,
1g,
1e,
0b,
1_,
1^,
1],
0[,
0Y,
1X,
0y/
0w/
1u/
1t/
1s/
1o/
0n/
0m/
0k/
1j/
0i/
1h/
1f/
1e/
0`/
1^/
1]/
1\/
0X/
0W/
1V/
1Q/
0O/
0N/
0M/
0I/
1H/
1G/
1E/
0D/
1C/
0B/
0@/
0?/
1:/
08/
07/
06/
12/
11/
00/
0u2
0n2
0l2
0k2
0j2
0i2
0g2
0e2
0b2
0^2
0W2
0V2
0U2
1T2
1O5
1L5
0K5
0J5
0I5
0F5
1C5
1A5
0=5
0;5
0:5
195
155
045
035
025
0/5
1.5
1-5
0,5
0#8
0z7
0x7
0w7
0v7
0u7
0s7
0q7
0n7
0j7
0c7
0b7
0a7
1`7
1;.
19.
18.
06.
15.
11.
1/.
0-.
1,.
0*.
0&.
0%.
0#.
0}-
0w-
0t-
0s-
1r-
0a.
0_.
0].
0V.
1U.
0T.
0S.
0Q.
0O.
1M.
1K.
1I.
0H.
0F.
1B.
1A.
0@.
0?.
1>.
1A+
1@+
1:+
04+
03+
1.+
0,+
1*+
1)+
0(+
1#+
1"+
0~*
1`+
1_+
1[+
1W+
1Q+
1P+
1O+
1I+
1H+
1D+
117
0.7
0-7
0+7
0*7
1)7
1(7
0$7
1#7
1"7
1~6
1}6
0|6
1{6
1z6
0y6
0x6
1w6
0u6
0t6
0r6
1n6
1[7
0Y7
1X7
1V7
1S7
1R7
0P7
1O7
1M7
0G7
0D7
1C7
1B7
1A7
1?7
1<7
1:7
087
174
144
124
014
104
1/4
1-4
1,4
0'4
0&4
0"4
1y3
0x3
1w3
1v3
0t3
1s3
1q3
0p3
0o3
1n3
0T4
0R4
0P4
0M4
0K4
1G4
1E4
1>4
0=4
0;4
191
071
161
051
021
011
101
0/1
0.1
1-1
1,1
0+1
1)1
1'1
0%1
1$1
1#1
0}0
0y0
0x0
1w0
1t0
0s0
0q0
1p0
1]1
0[1
1Y1
1W1
0U1
1S1
0Q1
0O1
0L1
0K1
1J1
1I1
1G1
1F1
0D1
1B1
1=1
0<1
0%:
1~9
1}9
0z9
1w9
0q9
0o9
1n9
0m9
0l9
0g9
1f9
0d9
1c9
1I:
0?:
19:
17:
15:
1/:
0+:
1*:
#45000
1"
1T!
b110111000001100011010001101010000111 N:
b1000110000011100000100010001100000 O:
b1000000111000000000101011001011111001101 P:
b10011000000111110000000100100000000000 Q:
b1000110100010011011011011011001000101001 R:
b1001110001111100000100110011100010000 S:
b1001110111011000110001000011111110111101 T:
b1000000111000000010100000000000000 U:
b111110100010011011011011011001000010000 V:
b101001111100000101010100110011100100 W:
b11010010010100101000000110011110000000 X:
b100101000001010101010001000000010000 Y:
b10101011100010011010111110010001000100100 "F
b1000100001000100101010000101010010000000 #F
b100000101010100001011011101111011011100110100 $F
b10101000100010101010100110000000100000000000 %F
b11101010000111001111100111110100110100100000 &F
b1000101000010000001000000000001000000000 'F
b10010110100111000101001101000011000000101101011100101101111011 P!
b1111101110000100011001101011110101010110011101101111111100100100 Q!
b10000100100001001101011000001001 H!
b10010000101010011010100100100 J!
b10110001111100000101011001100011 I!
b11000000100010010101111010000001 K!
1gY
1dY
1aY
1`Y
1_Y
1^Y
1]Y
1\Y
1[Y
1ZY
1XY
1WY
1UY
1TY
1SY
1PY
1OY
1MY
1KY
1IY
1GY
1FY
1EY
1DY
1BY
1@Y
1?Y
1<Y
1;Y
17Y
12Y
11Y
10Y
1.Y
1-Y
1,Y
1+Y
1*Y
1RJ
1FJ
1?J
1:J
18J
14J
1~I
1{I
1yI
1xI
1uI
1rI
1pI
0mI
1lI
1jI
1hI
0gI
1dI
0aI
0`I
0_I
0]I
0[I
1LI
1DI
1CI
1@I
1>I
1<I
1:I
18I
14I
10I
1.I
1,I
1dG
1bG
1aG
1^G
1]G
1\G
1ZG
1YG
1WG
1VG
1UG
1TG
1RG
1QG
1PG
1NG
1MG
1KG
1FG
1DG
0CG
1BG
0AG
1@G
0?G
0=G
0;G
1:G
09G
1/G
1,G
1*G
1(G
1#G
1!G
1}F
1zF
1vF
1qF
1mF
1\F
1YF
1UF
1QF
1NF
1MF
1LF
1KF
1JF
1HF
1FF
1EF
1BF
1>F
1=F
1<F
09F
18F
07F
16F
05F
1"D
0vC
1pC
1nC
1lC
1fC
0bC
1aC
0WC
1RC
1QC
0NC
1KC
0EC
0CC
1BC
0AC
0@C
0;C
1:C
08C
17C
10C
0.C
1-C
1+C
1(C
1'C
0%C
1$C
1"C
0zB
0wB
1vB
1uB
1tB
1rB
1oB
1mB
0kB
1aB
0^B
0]B
0[B
0ZB
1YB
1XB
0TB
1SB
1RB
1PB
1OB
0NB
1MB
1LB
0KB
0JB
1IB
0GB
0FB
0DB
1@B
0'@
0%@
0#@
0~?
0|?
1x?
1v?
1o?
0n?
0l?
1b?
1_?
1]?
0\?
1[?
1Z?
1X?
1W?
0R?
0Q?
0M?
1F?
0E?
1D?
1C?
0A?
1@?
1>?
0=?
0<?
1;?
14?
02?
10?
1.?
0,?
1*?
0(?
0&?
0#?
0"?
1!?
1~>
1|>
1{>
0y>
1w>
1r>
0q>
1h>
0f>
1e>
0d>
0a>
0`>
1_>
0^>
0]>
1\>
1[>
0Z>
1X>
1V>
0T>
1S>
1R>
0N>
0J>
0I>
1H>
1E>
0D>
0B>
1A>
0D<
0B<
0@<
09<
18<
07<
06<
04<
02<
10<
1.<
1,<
0+<
0)<
1%<
1$<
0#<
0"<
1!<
1z;
1x;
1w;
0u;
1t;
1p;
1n;
0l;
1k;
0i;
0e;
0d;
0b;
0^;
0X;
0U;
0T;
1S;
1K;
1J;
1F;
1B;
1<;
1;;
1:;
14;
13;
1/;
1&;
1%;
1}:
0w:
0v:
1q:
0o:
1m:
1l:
0k:
1f:
1e:
0c:
0jY
1NR
1MR
1HR
0CR
0AR
0@R
1?R
1;R
18R
16R
05R
11R
1/R
0-R
0,R
1A=
1@=
1?=
1:=
15=
13=
01=
1.=
1*=
1)=
1#=
1"=
1wR
1uR
1qR
1pR
1mR
0kR
1gR
0dR
0aR
1`R
1_R
1^R
1\R
1YR
1TR
0SR
1PR
02>
1(>
0&>
0$>
0">
1|=
1z=
0y=
1r=
0p=
1vS
0tS
1sS
0rS
0qS
0nS
1lS
1jS
1hS
0gS
1fS
0eS
0dS
1cS
0bS
1aS
0_S
0^S
0]S
1\S
1[S
0ZS
0WS
1SS
0RS
1QS
1OS
19A
16A
02A
10A
0/A
1.A
1-A
1,A
0+A
1)A
1(A
1$A
0#A
0"A
0}@
0y@
1w@
1t@
1s@
0q@
1p@
1AT
1>T
1<T
0;T
1:T
19T
17T
16T
15T
03T
10T
0.T
1(T
0&T
1%T
0$T
1#T
1"T
0~S
1|S
1{S
0yS
1xS
0%B
0~A
0|A
1vA
1oA
0nA
0lA
1BU
1AU
0@U
1?U
1>U
0;U
18U
07U
06U
13U
02U
00U
1/U
1-U
1,U
1(U
1'U
0$U
0#U
0!U
1~T
1}T
1#E
0~D
0}D
1yD
1xD
1wD
0tD
1sD
1oD
0nD
1mD
1lD
0kD
1iD
0gD
0fD
0aD
1`D
0iU
1fU
1dU
1cU
0`U
1]U
0\U
0WU
0VU
0UU
0SU
0MU
1JU
1IU
0HU
0GU
0jE
1dE
1bE
1`E
1ZE
1EH
1BH
1?H
1>H
1=H
1<H
1;H
1:H
18H
14H
13H
12H
10H
1/H
1-H
1,H
1*H
1)H
1(H
1%H
1$H
0#H
0"H
1!H
0~G
1}G
0|G
1{G
0zG
1yG
0xG
1wG
0vG
0tG
0rG
1qG
0pG
1qH
1nH
1mH
1lH
1jH
1hH
1fH
1eH
1bH
1^H
1]H
1ZH
1VH
15K
10K
1,K
1*K
1)K
0%K
1$K
0#K
1"K
0!K
1|J
0{J
1zJ
1xJ
1vJ
0uJ
1tJ
0sJ
0pJ
0mJ
1dK
1bK
1^K
1\K
1ZK
1XK
1TK
1NK
1LK
1TD
0QD
0PD
1LD
1KD
1JD
0GD
1FD
1BD
0AD
1@D
1?D
0>D
1<D
0:D
09D
04D
13D
1<V
1;V
0:V
19V
18V
17V
05V
04V
10V
1.V
1-V
0,V
1+V
1)V
1'V
0&V
0%V
1$V
0#V
1"V
0|U
1{U
1xU
1wU
1vU
1uU
0tU
0sU
0#E
0wD
0sD
1pD
0oD
0mD
0lD
1hD
1aD
0_D
1g@
1d@
0`@
1^@
0]@
1\@
1[@
1Z@
0Y@
1W@
1V@
1R@
0Q@
0P@
0M@
0I@
1G@
1D@
1C@
0A@
1@@
1vT
0tT
1sT
0rT
0qT
1pT
1nT
1mT
0lT
0kT
0iT
1gT
0cT
0aT
1^T
1\T
1[T
1ZT
1UT
1TT
1MT
1LT
0JT
1IT
09A
06A
14A
01A
1/A
0-A
1+A
0(A
0$A
1~@
0t@
0s@
1r@
0p@
1s<
1r<
1q<
1l<
1g<
1e<
0c<
1`<
1\<
1[<
1U<
1T<
1FS
1ES
0DS
1BS
1@S
1>S
0=S
1;S
0:S
09S
17S
04S
13S
11S
00S
1,S
1+S
1'S
0&S
1%S
1$S
1!S
0~R
1{R
0A=
0@=
03=
0.=
1+=
0)=
0"=
0~<
0s<
0r<
0e<
0`<
1]<
0[<
0T<
0R<
1l=
1i=
1h=
1f=
0c=
1a=
1`=
0[=
0Z=
0Y=
0X=
1W=
0V=
0T=
0S=
1R=
1Q=
0K=
0J=
1G=
0F=
1C=
18>
11>
0->
1*>
1&>
1%>
1!>
1~=
0}=
0|=
1x=
1v=
1u=
0r=
0g@
0d@
1b@
0_@
1]@
0[@
1Y@
0V@
0R@
1N@
0D@
0C@
1B@
0@@
1hA
1gA
0fA
1eA
0cA
1bA
0_A
0\A
1ZA
0WA
0VA
1UA
0SA
0RA
1QA
1NA
1LA
1IA
0FA
0DA
1CA
1AA
1@A
1?A
1>A
0<A
1;A
10B
0.B
1-B
1(B
1'B
0&B
1$B
1#B
0"B
0xA
1uA
1sA
0pA
0TD
0JD
0FD
1CD
0BD
0@D
0?D
1;D
14D
02D
1PE
1OE
1ME
1LE
1JE
0IE
0HE
1FE
0EE
0BE
0?E
1=E
0<E
17E
04E
03E
12E
11E
0,E
1+E
0*E
0)E
0vE
1tE
1qE
1pE
1nE
1lE
1kE
1hE
1fE
0dE
0cE
0^E
0ZE
1YE
1UE
0NE
1DE
0@E
0=E
1<E
0:E
09E
05E
0.E
1,E
0pE
1iE
0hE
1aE
1ZE
0XE
0gA
0dA
0bA
1_A
1]A
0[A
0YA
1VA
1RA
0NA
1DA
0CA
0BA
0@A
13B
00B
1*B
0'B
0#B
1}A
0sA
1qA
1k=
0j=
1]=
1X=
1U=
1S=
0L=
1J=
08>
0*>
0%>
0~=
0u=
#46800
b110101110010111101100001101 d
b1000110110111111001100110001101 e
0"
0(Y
1'Y
1&Y
0$Y
0#Y
1"Y
1!Y
0~X
0}X
1|X
0yX
1xX
1wX
1vX
1uX
1tX
0rX
0oX
1nX
1mX
0kX
0jX
1iX
0hX
0t!
1s!
1r!
0p!
0o!
1n!
1m!
0l!
0k!
1j!
0g!
1f!
1e!
1d!
1c!
1b!
0`!
0]!
1\!
1[!
0Y!
0X!
1W!
0V!
1eX
1_X
0]X
1\X
1ZX
0XX
1WX
0UX
1TX
1SX
1RX
1NX
0HX
0F!
0C!
0A!
09!
07!
16!
03!
02!
00!
1/!
1-!
1,!
0(!
0#!
0~
1}
1|
1v
0u
0t
1r
1q
0p
1o
0k
0h
0T!
0q(
1p(
1o(
0m(
0l(
1k(
1j(
0i(
0h(
1g(
0d(
1c(
1b(
1a(
1`(
1_(
0](
0Z(
1Y(
1X(
0V(
0U(
1T(
0S(
15"
1/"
0-"
1,"
1*"
0("
1'"
0%"
1$"
1#"
1""
1|!
0v!
b0 yQ
b1 pQ
b1 gQ
b0 aQ
b1 [Q
1MQ
0PQ
1SQ
0YQ
1_Q
1eQ
0nQ
1tQ
b1000110110111111001100110001101 KQ
b110111001001000000110011001110010 NQ
b1000110110111111001100110001101 QQ
b110111001001000000110011001110010 WQ
b110111001001000000110011001110010 ZQ
b0 ]Q
b10001101101111110011001100011010 `Q
b1000110110111111001100110001101 cQ
b101110010010000001100110011100101 fQ
b110111001001000000110011001110010 lQ
b110111001001000000110011001110010 oQ
b10001101101111110011001100011010 rQ
b0 xQ
1%)
0$)
1#)
0!)
1}(
1{(
0x(
1v(
0q'
0n'
0m'
0l'
0i'
0h'
0e'
0c'
0a'
0`'
0_'
0^'
0]'
0W'
0V'
0U'
0R'
0/'
1,'
1+'
0*'
0)'
1''
0%'
1"'
0!'
1}&
1|&
1{&
1z&
0w&
1s&
1r&
0q&
0p&
0m&
0l&
1h&
0`&
1_&
0X&
0V&
0U&
1Q&
0K&
1J&
0H&
1E&
0C&
1A&
0?&
1>&
0;&
0:&
09&
08&
07&
16&
13&
01&
1.&
1+&
0f%
1e%
1`%
0^%
1\%
0[%
1X%
0S%
0R%
0P%
0O%
1N%
1I%
0H%
0E%
1D%
1C%
0A%
0@%
1?%
1>%
0=%
0<%
1;%
08%
17%
16%
15%
14%
13%
01%
0.%
1-%
1,%
0*%
0)%
1(%
0'%
0&%
1$%
0#%
0|$
1z$
0x$
1w$
0t$
1o$
1n$
1l$
1k$
0j$
0e$
1d$
0b$
0a$
0]$
0\$
0Y$
0X$
0V$
0T$
0N$
0M$
0L$
0K$
0J$
0F$
0E$
0C$
0B$
0?$
1=$
1<$
0:$
18$
06$
13$
02$
0+$
0*$
0($
1&$
1%$
0#$
1"$
0~#
1}#
0{#
1x#
0v#
1t#
0r#
1q#
0n#
0m#
0l#
0k#
0j#
1i#
1f#
0d#
1a#
1^#
0;#
1:#
19#
07#
06#
15#
14#
03#
02#
11#
0.#
1-#
1,#
1+#
1*#
1)#
0'#
0$#
1##
1"#
0~"
0}"
1|"
0{"
0z"
0y"
1x"
0v"
1s"
0q"
1o"
0m"
1l"
0i"
0h"
0g"
0f"
0e"
1d"
1a"
0_"
1\"
1Y"
0W"
1V"
1U"
0S"
0R"
1Q"
1P"
0O"
0N"
1M"
0J"
1I"
1H"
1G"
1F"
1E"
0C"
0@"
1?"
1>"
0<"
0;"
1:"
09"
08"
1>(
0B(
1F(
1L(
0R(
0m8
1w2
0)/
1'/
1&/
0$/
1"/
0~.
1{.
0z.
0s.
0r.
0p.
1n.
1m.
0k.
1j.
1v/
0u/
0p/
1n/
0l/
1k/
0h/
1c/
1b/
1`/
1_/
0^/
0Y/
1X/
0N2
1M2
1H2
0F2
1D2
0C2
1@2
0;2
0:2
082
072
162
112
002
0M5
1I5
0A5
1@5
095
075
065
125
0G8
0D8
0C8
0B8
0?8
0>8
0;8
098
078
068
058
048
038
0-8
0,8
0+8
0(8
1u5
0s5
1p5
1o5
0n5
0m5
1k5
0i5
1f5
0e5
1c5
1b5
1a5
1`5
0]5
1Y5
1X5
0W5
0V5
0S5
1R5
0'5
1&5
0$5
1!5
0}4
1{4
0y4
1x4
0u4
0t4
0s4
0r4
0q4
1p4
1m4
0k4
1h4
1e4
0d4
0+2
0(2
1'2
1&2
0$2
0#2
1"2
1!2
0~1
0}1
1|1
0y1
1x1
1w1
1v1
1u1
1t1
0r1
0o1
1n1
1m1
0k1
0j1
1i1
0h1
0g1
1f1
1S/
0Q/
0P/
0L/
0K/
0H/
0G/
0E/
0C/
0=/
0</
0;/
0:/
09/
05/
04/
02/
01/
10/
0y,
1x,
0v,
1s,
0q,
1o,
0m,
1l,
0i,
0h,
0g,
0f,
0e,
1d,
1a,
0_,
1\,
1Y,
0X,
0,,
1+,
1*,
0(,
0',
1&,
1%,
0$,
0#,
1",
0}+
1|+
1{+
1z+
1y+
1x+
0v+
0s+
1r+
1q+
0o+
0n+
1m+
0l+
0k+
1j+
01*
10*
0.*
1+*
0)*
1'*
0%*
1$*
0!*
0~)
0})
0|)
0{)
1z)
1w)
0u)
1r)
1o)
0n)
0l)
1k)
1j)
0h)
0g)
1f)
1e)
0d)
0c)
1b)
0_)
1^)
1])
1\)
1[)
1Z)
0X)
0U)
1T)
1S)
0Q)
0P)
1O)
0N)
0M)
0L)
0K)
1J)
0@+
1;+
0:+
08+
06+
05+
01+
10+
1-+
1++
0*+
0)+
1(+
1$+
0#+
0!+
1~*
1b+
0`+
0_+
1^+
1]+
0[+
1Z+
1Y+
0W+
1V+
1U+
0Q+
0P+
0O+
1N+
1K+
0I+
0H+
1G+
0D+
08.
17.
16.
05.
03.
01.
10.
1..
1-.
1*.
0'.
1&.
1%.
1#.
1".
1}-
0z-
1x-
1w-
1s-
0r-
1Y.
0X.
0U.
1P.
1O.
0M.
0L.
0K.
0J.
0I.
1H.
0B.
0A.
1@.
137
127
107
1/7
0,7
1*7
0&7
1$7
0#7
0~6
0z6
1x6
0s6
1r6
0m6
1l6
0[7
0X7
0W7
1U7
1T7
0R7
1N7
0M7
0I7
1F7
1D7
0B7
0A7
1>7
1=7
0:7
171
041
131
111
1/1
1.1
0,1
1+1
0*1
0$1
1|0
0{0
1x0
0t0
0]1
1Z1
0Y1
0X1
0W1
0T1
0S1
1R1
0P1
0I1
0H1
0F1
1D1
1C1
0B1
0A1
0=1
1<1
074
044
114
004
0/4
0.4
0-4
0+4
1(4
1&4
0%4
1#4
1"4
0~3
1}3
1|3
1{3
1x3
0w3
0v3
0u3
1t3
1[4
1V4
1U4
0O4
1M4
1L4
0G4
0F4
0E4
1?4
0>4
0~9
0}9
0|9
1y9
0x9
1u9
1s9
1q9
0p9
1o9
0n9
1m9
1g9
0f9
1e9
1b9
0I:
0A:
0=:
0;:
09:
07:
05:
0/:
0-:
0*:
#48600
1"
1T!
b111010100010010111100000000001000101 N:
b1000100100000011001100110001000 O:
b100011101010011011001111111101010110101 P:
b10100000001000000110000000010000000000 Q:
b1000010110001011010011010101111101001101 R:
b10001001100100100000001000000010000000 S:
b1001111000111111011100101010100001110100 T:
b100000000000011000100011000010000 U:
b1011111000011001010010110011100001111100 V:
b1111100110100001001100011110000000 W:
b11110101010101010101010101010000000000 X:
b0 Y:
b110011010000011110101100011011100001111011 "F
b101010100001000010100100010100000000 #F
b1001101001000110011011110111010100111100001001 $F
b10100111000100100001000101001000001000000 %F
b10011000011000011001100001011010001111011000 &F
b1000110100011100010010110100100100000000000 'F
b10000010101010100110011101101101110001011111100100100 xK
b10001001100010011010101110010000000000000 yK
b1111101101001011111011001010000110100010000100000000000 zK
b10100000100010101010001010000000000000000000 {K
b111011100100101110100000001001101000001101000101100101001 P!
b10010110100111000101001101000011000000101101011100101101111011 Q!
b1111101110000100011001101011110101010110011101101111111100100100 R!
b110101110010111101100001101 H!
b10000100100001001101011000001001 J!
b10010000101010011010100100100 L!
b1000110110111111001100110001101 I!
b10110001111100000101011001100011 K!
b11000000100010010101111010000001 M!
1iY
1hY
0gY
1fY
1eY
1cY
0_Y
0]Y
0\Y
1YY
0XY
0SY
1RY
0PY
0OY
0MY
1JY
0IY
0GY
0FY
0DY
1CY
0@Y
1=Y
0<Y
0;Y
19Y
18Y
14Y
00Y
1/Y
0.Y
0-Y
0+Y
0*Y
1DN
1BN
1>N
1<N
1:N
18N
14N
1.N
1,N
1kM
1fM
1bM
1`M
1_M
0[M
1ZM
0YM
1XM
0WM
1TM
0SM
1RM
1PM
1NM
0MM
1LM
0KM
0HM
0EM
11M
1.M
1-M
1,M
1*M
1(M
1&M
1%M
1"M
1|L
1{L
1xL
1tL
1[L
1XL
1UL
1TL
1SL
1RL
1QL
1PL
1NL
1JL
1IL
1HL
1FL
1EL
1CL
1BL
1@L
1?L
1>L
1;L
1:L
09L
08L
17L
06L
15L
04L
13L
02L
11L
00L
1/L
0.L
0,L
0*L
1)L
0(L
0RJ
1PJ
1MJ
1JJ
1HJ
1GJ
0FJ
1EJ
1BJ
0?J
1>J
1=J
1<J
0:J
16J
15J
04J
11J
1"J
1!J
0~I
1}I
1|I
1zI
0yI
0xI
1vI
0uI
1tI
0rI
0pI
0oI
0jI
0iI
1gI
0eI
0dI
0cI
1bI
1aI
0^I
1[I
0ZI
0YI
1QI
0LI
1KI
1HI
1FI
0DI
0CI
1BI
0@I
0>I
1=I
0<I
08I
16I
15I
11I
00I
1/I
0.I
0,I
1fG
0dG
1cG
0bG
0aG
1[G
0ZG
0YG
1XG
0WG
0UG
1SG
0QG
1OG
1JG
1GG
0DG
0@G
1?G
1=G
1<G
0:G
19G
0/G
1.G
0*G
1%G
0!G
0}F
1|F
0zF
1wF
0vF
1uF
1sF
0mF
1^F
1]F
0\F
1[F
1ZF
1XF
0UF
1SF
1RF
1OF
0MF
0LF
0KF
1IF
0HF
1GF
0FF
1DF
1CF
0>F
0=F
19F
08F
15F
0"D
0xC
0tC
0rC
0pC
0nC
0lC
0fC
0dC
0aC
0RC
0QC
0PC
1MC
0LC
1IC
1GC
1EC
0DC
1CC
0BC
1AC
1;C
0:C
19C
16C
00C
0-C
0,C
1*C
1)C
0'C
1#C
0"C
0|B
1yB
1wB
0uB
0tB
1qB
1pB
0mB
1cB
1bB
1`B
1_B
0\B
1ZB
0VB
1TB
0SB
0PB
0LB
1JB
0EB
1DB
0?B
1>B
1.@
1)@
1(@
0"@
1~?
1}?
0x?
0w?
0v?
1p?
0o?
0b?
0_?
1\?
0[?
0Z?
0Y?
0X?
0V?
1S?
1Q?
0P?
1N?
1M?
0K?
1J?
1I?
1H?
1E?
0D?
0C?
0B?
1A?
04?
11?
00?
0/?
0.?
0+?
0*?
1)?
0'?
0~>
0}>
0{>
1y>
1x>
0w>
0v>
0r>
1q>
1f>
0c>
1b>
1`>
1^>
1]>
0[>
1Z>
0Y>
0S>
1M>
0L>
1I>
0E>
1<<
0;<
08<
13<
12<
00<
0/<
0.<
0-<
0,<
1+<
0%<
0$<
1#<
0w;
1v;
1u;
0t;
0r;
0p;
1o;
1m;
1l;
1i;
0f;
1e;
1d;
1b;
1a;
1^;
0[;
1Y;
1X;
1T;
0S;
1M;
0K;
0J;
1I;
1H;
0F;
1E;
1D;
0B;
1A;
1@;
0<;
0;;
0:;
19;
16;
04;
03;
12;
0/;
0%;
1~:
0}:
0{:
0y:
0x:
0t:
1s:
1p:
1n:
0m:
0l:
1k:
1g:
0f:
0d:
1c:
0MR
1JR
1FR
1AR
0?R
1:R
09R
15R
13R
0/R
0.R
1-R
1,R
1;=
0:=
06=
05=
12=
11=
10=
1.=
1-=
0+=
0*=
1)=
1(=
0#=
1~<
1|<
0tR
1sR
1rR
0qR
0oR
0mR
1kR
1jR
1iR
1hR
1fR
1aR
0`R
0]R
0\R
0XR
1VR
0TR
1SR
0QR
0PR
1,>
0+>
0(>
1#>
1">
0z=
1y=
1q=
1tS
1pS
1mS
0iS
0fS
1dS
0aS
1]S
0\S
0[S
1XS
1VS
0US
0SS
0QS
1PS
17A
04A
13A
11A
1-A
0,A
0+A
0*A
0)A
1$A
1}@
1|@
0{@
1x@
1t@
0r@
1p@
0AT
0>T
0<T
1;T
0:T
09T
08T
06T
05T
02T
0/T
1.T
1,T
0*T
1)T
1&T
1$T
0#T
0"T
0!T
1}S
1.B
1)B
1~A
0oA
1CU
1@U
0>U
1;U
0:U
19U
16U
05U
03U
0-U
0,U
1+U
0*U
1)U
0(U
1!U
0}T
1|T
1%E
1"E
0xD
0vD
1sD
0pD
1oD
1mD
0jD
0hD
1gD
1dD
0`D
1_D
1^D
0fU
0dU
0cU
0bU
1_U
1[U
0ZU
1YU
0XU
1WU
1UU
1SU
0RU
1MU
1KU
0JU
1HU
1GU
0tE
0lE
0fE
0`E
0UE
1GH
1FH
0EH
1DH
1CH
1AH
0=H
08H
16H
03H
11H
0-H
0,H
0*H
0)H
1&H
0%H
1#H
1"H
0!H
1~G
0}G
1|G
0{G
0wG
1vG
1tG
1sG
0qG
1pG
1sH
0qH
1oH
0mH
0hH
0fH
1dH
1cH
1`H
0]H
1\H
1:K
05K
14K
12K
00K
1.K
1-K
1+K
0*K
1(K
1&K
1%K
0$K
1#K
0"K
1!K
1~J
0zJ
0xJ
1uJ
1sJ
1rJ
0nJ
1mJ
0lJ
0jJ
0iJ
0hJ
1hK
1fK
0dK
0bK
0^K
1]K
0\K
0XK
1UK
1QK
0NK
0LK
1EK
1AK
1"W
1}V
1zV
1yV
1xV
1wV
1vV
1uV
1tV
1sV
1qV
1pV
1nV
1jV
1iV
1gV
1dV
1cV
1aV
1_V
0^V
1\V
0[V
1ZV
1XV
0WV
1VV
0UV
1TV
0SV
0QV
0OV
1NV
0MV
1EQ
1BQ
1?Q
1>Q
1=Q
1<Q
1;Q
1:Q
18Q
14Q
13Q
12Q
10Q
1/Q
1-Q
1,Q
1*Q
1)Q
1(Q
1%Q
1$Q
0#Q
1"Q
1!Q
1~P
1}P
1{P
1zP
1yP
1xP
1wP
1vP
1tP
1rP
1qP
1PW
1KW
1DW
1AW
0@W
0>W
0<W
1;W
19W
08W
15W
13W
02W
00W
1/W
0-W
0*W
1fO
1dO
1`O
1bP
1_P
1\P
1[P
1ZP
1YP
1XP
1WP
1UP
1QP
1PP
1OP
1MP
1LP
1JP
1IP
1GP
1FP
1EP
1BP
1AP
0@P
1?P
1>P
1=P
1<P
1:P
19P
18P
17P
16P
15P
13P
11P
10P
1DX
1AX
1>X
1=X
1<X
1;X
1:X
19X
18X
17X
15X
14X
1.X
1+X
1(X
1'X
1&X
1%X
0}W
0{W
0zW
0wW
0vW
0rW
0qW
0mW
0jW
0EQ
0BQ
0?Q
0>Q
0=Q
0<Q
0;Q
0:Q
08Q
0/Q
1.Q
0,Q
0)Q
0$Q
0!Q
0~P
0}P
0zP
0yP
0xP
0vP
0tP
0rP
0qP
1VD
1SD
0KD
0ID
1FD
0CD
1BD
1@D
0=D
0;D
1:D
17D
03D
12D
11D
1=V
1:V
08V
15V
13V
12V
01V
1/V
0)V
0(V
0$V
0"V
0!V
1~U
1tU
1sU
0%E
0"E
1zD
0yD
0sD
1kD
1jD
0_D
0^D
1e@
0b@
1a@
1_@
1[@
0Z@
0Y@
0X@
0W@
1R@
1M@
1L@
0K@
1H@
1D@
0B@
1@@
1tT
1kT
0jT
1hT
0gT
1fT
0eT
0^T
0\T
0YT
0VT
0RT
1NT
07A
03A
00A
1)A
0'A
0$A
0~@
0}@
1y@
0v@
0t@
1m<
0l<
0h<
0g<
1d<
1c<
1b<
1`<
1_<
0]<
0\<
1[<
1Z<
0U<
1R<
1P<
0ES
0BS
0AS
0@S
1?S
0<S
1:S
19S
18S
06S
15S
03S
02S
01S
0.S
0+S
0*S
1)S
0'S
1&S
0$S
0#S
0!S
1~R
0|R
0{R
1==
14=
02=
0(=
1&=
1"=
0!=
0~<
1o<
1f<
0d<
0Z<
1X<
1T<
0S<
0R<
0k=
0h=
0g=
0f=
1d=
1b=
1^=
1Z=
1Y=
0U=
0S=
0R=
0Q=
0P=
1O=
1L=
1I=
0H=
0G=
1F=
0D=
0C=
12>
01>
0/>
0,>
1(>
0&>
0!>
1~=
1}=
0x=
0t=
1s=
0q=
1o=
0e@
0a@
0^@
1W@
0U@
0R@
0N@
0M@
1I@
0F@
0D@
1fA
0eA
1bA
1aA
0_A
0]A
1\A
1[A
0RA
0PA
1NA
0MA
0LA
1BA
16B
03B
10B
0-B
0*B
0)B
1#B
1|A
1{A
0zA
0qA
1oA
0VD
0SD
1MD
0LD
0FD
1>D
1=D
02D
01D
1QE
0PE
1NE
0ME
0LE
1IE
1GE
0FE
1@E
1:E
08E
07E
16E
01E
1-E
0,E
0+E
1*E
1)E
1|E
1yE
1rE
0qE
0iE
0bE
0aE
1`E
1]E
0YE
1XE
1WE
0bP
0_P
0\P
0[P
0ZP
0YP
0XP
0WP
0UP
0LP
1KP
0IP
0FP
0AP
0>P
0=P
0<P
09P
08P
07P
05P
03P
01P
00P
1AO
1@O
1>O
1=O
1;O
14O
13O
12O
11O
1/O
1.O
1-O
1*O
1'O
1"O
1~N
1}N
1|N
0{N
0yN
0wN
0vN
0uN
0rN
0qN
0nN
0mN
0lN
0jN
0gN
1zO
1yO
1xO
1wO
1vO
1uO
1kO
1hO
1eO
1cO
0^O
1]O
1\O
1[O
1ZO
1XO
1WO
1VO
1TO
1SO
1PO
1OO
1NO
0@O
0=O
1:O
19O
18O
17O
16O
15O
03O
0*O
1)O
0'O
1$O
0}N
0zN
1yN
0xN
1uN
0tN
0sN
1qN
0oN
1mN
1lN
0zO
0yO
0xO
0wO
0vO
0uO
0dO
0[O
0WO
0SO
0OO
0NO
1PE
1ME
0GE
1FE
0@E
18E
17E
1,E
1+E
0|E
0yE
1sE
0rE
0XE
0WE
1eA
0aA
0^A
1WA
0UA
1RA
0NA
1MA
0IA
1FA
0DA
06B
0#B
0|A
1xA
0uA
1g=
0^=
0\=
1R=
1P=
0L=
1K=
0J=
1+>
0}=
1w=
0v=
#50400
b10110010110000101000010001100101 d
b10001001001101110101001000010010 e
0"
0)Y
1(Y
0'Y
0&Y
1%Y
0"Y
0!Y
1~X
0|X
1yX
0xX
0tX
1rX
0qX
0pX
1oX
0nX
0mX
1lX
0iX
1hX
0u!
1t!
0s!
0r!
1q!
0n!
0m!
1l!
0j!
1g!
0f!
0b!
1`!
0_!
0^!
1]!
0\!
0[!
1Z!
0W!
1V!
0dX
1bX
1aX
0_X
0^X
1]X
0\X
0[X
0ZX
0YX
1XX
0WX
1VX
0TX
0SX
0RX
1QX
0MX
1KX
1JX
1HX
0G!
1F!
1C!
0B!
0>!
1:!
06!
05!
14!
11!
10!
0/!
1.!
1+!
1%!
1$!
1#!
1"!
0{
0y
1x
1w
1t
0r
1l
1h
0T!
0r(
1q(
0p(
0o(
1n(
0k(
0j(
1i(
0g(
1d(
0c(
0_(
1](
0\(
0[(
1Z(
0Y(
0X(
1W(
0T(
1S(
04"
12"
11"
0/"
0."
1-"
0,"
0+"
0*"
0)"
1("
0'"
1&"
0$"
0#"
0""
1!"
0{!
1y!
1x!
1v!
b1 yQ
b1 vQ
b0 gQ
b1 dQ
b1 aQ
b0 [Q
b0 XQ
b0 OQ
b1 RQ
0MQ
0VQ
1YQ
1nQ
1qQ
0tQ
b110001001001101110101001000010010 KQ
b110001001001101110101001000010010 NQ
b11101101100100010101101111011011 QQ
b100010010011011101010010000100100 TQ
b0 WQ
b110001001001101110101001000010010 ZQ
b11101101100100010101101111011011 `Q
b1110110110010001010110111101101 cQ
b110001001001101110101001000010010 fQ
b1110110110010001010110111101101 lQ
b1110110110010001010110111101101 oQ
b110001001001101110101001000010010 rQ
b1110110110010001010110111101101 uQ
b1110110110010001010110111101101 xQ
0%)
0")
1!)
1x(
1w(
0v(
1q'
1o'
1n'
1l'
1k'
1j'
1i'
1g'
1f'
1d'
1b'
1^'
1['
1Z'
1X'
1W'
1U'
1T'
1S'
1P'
1N'
1M'
1K'
1J'
1I'
1H'
1F'
1E'
1C'
1A'
1='
1:'
19'
17'
16'
14'
13'
12'
0,'
0''
0"'
1!'
0z&
0v&
0s&
1m&
1l&
0k&
1j&
1i&
0h&
1e&
1d&
0c&
1a&
0^&
1]&
1Y&
0W&
1V&
1U&
0T&
1S&
1R&
0Q&
1N&
0M&
0L&
1K&
0J&
1I&
1H&
0G&
1D&
1C&
0B&
1@&
0=&
1<&
18&
06&
15&
14&
03&
12&
11&
00&
1-&
0,&
0+&
0g%
1f%
0e%
1c%
0b%
0a%
0`%
1^%
0]%
0\%
1[%
0X%
1W%
1V%
1U%
1S%
1R%
0Q%
1O%
0N%
1L%
0K%
0J%
0I%
1H%
1A%
1@%
1<%
0:%
19%
06%
05%
04%
02%
1*%
1)%
1%%
1}$
1|$
1x$
0v$
1u$
0r$
0q$
0p$
0n$
1f$
1e$
0<$
0;$
07$
15$
04$
11$
10$
1/$
1-$
0%$
0$$
0}#
0z#
0y#
0x#
0u#
0t#
0q#
0p#
0i#
0f#
0c#
0b#
0a#
0_#
0^#
1[#
1X#
1S#
1P#
1N#
1L#
1K#
1J#
1H#
1G#
1D#
1A#
1=#
1;#
0:#
18#
16#
13#
1.#
0-#
0+#
0*#
0)#
0&#
1$#
0##
1!#
1}"
1{"
0t"
0s"
0o"
1m"
0l"
1i"
1h"
1g"
1e"
0]"
0\"
0X"
1W"
0V"
0U"
1T"
0Q"
0P"
1O"
0M"
1J"
0I"
0E"
1C"
0B"
0A"
1@"
0?"
0>"
1="
0:"
19"
18"
18(
06(
0<(
0>(
1B(
1D(
0F(
1P(
1R(
1m8
0w2
0S/
0,*
0+*
0'*
1%*
0$*
1!*
1~)
1})
1{)
0s)
0r)
0/,
1,,
0+,
1),
1',
1$,
1}+
0|+
0z+
0y+
0x+
0u+
1s+
0r+
1p+
1n+
1l+
0-/
0&/
0%/
0!/
1}.
0|.
1y.
1x.
1w.
1u.
0m.
0l.
1w/
1q/
1p/
1l/
0j/
1i/
0f/
0e/
0d/
0b/
1Z/
1Y/
1+2
1$2
1#2
1}1
0{1
1z1
0w1
0v1
0u1
0s1
1k1
1j1
1Q2
0O2
1N2
0M2
1K2
0J2
0I2
0H2
1F2
0E2
0D2
1C2
0@2
1?2
1>2
1=2
1;2
1:2
092
172
062
142
032
022
012
102
1#8
1!8
1~7
1|7
1{7
1z7
1y7
1w7
1v7
1t7
1r7
1n7
1k7
1j7
1h7
1g7
1e7
1d7
1c7
1I8
1G8
1E8
1D8
1B8
1A8
1@8
1?8
1=8
1<8
1:8
188
148
118
108
1.8
1-8
1+8
1*8
1)8
0p5
0k5
0f5
1e5
0`5
0\5
0Y5
1S5
0R5
1M5
0L5
1K5
1J5
0I5
1F5
1E5
0D5
1B5
0?5
1>5
1:5
085
175
165
055
145
135
025
1/5
0.5
0-5
1,5
1'5
0&5
1%5
1$5
0#5
1~4
1}4
0|4
1z4
0w4
1v4
1r4
0p4
1o4
1n4
0m4
1l4
1k4
0j4
1g4
0f4
0e4
1d4
0x,
0u,
0t,
0s,
0p,
0o,
0l,
0k,
0d,
0a,
0^,
0],
0\,
0Z,
0Y,
1X,
1U,
1Q,
1N,
1I,
1F,
1D,
1B,
1A,
1@,
1>,
1=,
1:,
17,
13,
02,
0m)
1l)
0k)
0j)
1i)
0f)
0e)
1d)
0b)
1_)
0^)
0Z)
1X)
0W)
0V)
1U)
0T)
0S)
1R)
0O)
1N)
1M)
1L)
1K)
0J)
037
027
1.7
1-7
1+7
0)7
1'7
1&7
0%7
0$7
1#7
1!7
1~6
0{6
1z6
1v6
1u6
1t6
0r6
0o6
0n6
1m6
0l6
1[7
1Y7
0U7
1Q7
0O7
1L7
0K7
1E7
0D7
1B7
0@7
0>7
187
0;.
09.
18.
07.
04.
13.
02.
11.
0/.
0-.
0,.
1(.
0%.
1$.
0#.
0".
0{-
1z-
0y-
0w-
1v-
1u-
0s-
1r-
1a.
1].
1Z.
0Y.
1U.
0P.
0O.
1M.
1J.
1I.
0H.
1F.
1C.
0@.
0>.
0A+
1@+
0?+
1>+
1=+
18+
16+
15+
0/+
0-+
1,+
1*+
1)+
0(+
1'+
1&+
1!+
0~*
0}*
0|*
0b+
0^+
0]+
0Z+
0Y+
1W+
0V+
1S+
1Q+
0N+
0K+
0G+
1D+
1C+
091
071
031
121
011
1,1
0+1
1*1
1(1
0'1
0#1
1"1
0!1
0~0
0|0
1y0
0x0
1t0
1s0
1[1
0Z1
1S1
0R1
1O1
1M1
1K1
0J1
0C1
174
054
024
014
104
1.4
1-4
0,4
1+4
0*4
1'4
1%4
0"4
0}3
0|3
0{3
0y3
0x3
1w3
1u3
0t3
0s3
0r3
1]4
0[4
1Z4
1W4
0V4
0U4
1R4
0Q4
0M4
0L4
1J4
1G4
1F4
1C4
1@4
0?4
1<4
1#:
1":
1!:
1}9
1z9
1x9
0w9
1r9
1p9
1n9
0m9
1l9
0k9
0i9
1h9
1f9
1d9
0c9
1K:
1I:
1F:
1D:
1C:
1A:
1?:
1>:
1<:
15:
13:
12:
11:
1/:
1-:
1+:
#52200
1"
1T!
b110101101111010100001101001011010 N:
b11000000000000101010100000000000000 O:
b1001101010010000101011110010110100101000 P:
b100100110010000000100001001000100 Q:
b1001110101000000100010111011111010001000 R:
b10001000100100010101000100000001000000 S:
b1001000101001000010101111001011010010001 T:
b100010010011001000000010000100100100 U:
b100110011111010011111001110110111110000 V:
b10001101001101100000101001011010010100 W:
b11101111100010111111010011110101110000 X:
b10101011101000000101101011010010100 Y:
b100101000110100001111001011110100101001 "F
b10001000101000010110000100100000010000000 #F
b1001101100010100001010110101110111000101001101 $F
b10000101010010110001000100000101000000000 %F
b11111100001000111011100001011010011101111100 &F
b10110010000000000100100001000000000000 'F
b100110100100101011101010000001111010100011101101111011 xK
b10001010101011110000101011000100000000000 yK
b1010101111111010011110101101101111000101000001000000 zK
b1000100000000000100110000100100000000101000000000000000 {K
b1111101101110011000100010010101010000100011101101111111100100100 HQ
b1000101010101100100101101001000000000000000000000000 IQ
b10001111010110111000110111110001011110110010001010100100011010 P!
b111011100100101110100000001001101000001101000101100101001 Q!
b10010110100111000101001101000011000000101101011100101101111011 R!
b1111101110000100011001101011110101010110011101101111111100100100 S!
b10110010110000101000010001100101 H!
b110101110010111101100001101 J!
b10000100100001001101011000001001 L!
b10010000101010011010100100100 N!
b10001001001101110101001000010010 I!
b1000110110111111001100110001101 K!
b10110001111100000101011001100011 M!
b11000000100010010101111010000001 O!
0hY
0eY
0cY
0[Y
0YY
1XY
0UY
0TY
0RY
1QY
1OY
1NY
0JY
0EY
0BY
1AY
1@Y
1:Y
09Y
08Y
16Y
15Y
04Y
13Y
0/Y
0,Y
1a
1^
1[
1Z
1Y
1X
1W
1V
1U
1T
1R
1Q
1O
1N
1M
1J
1I
1G
1E
1C
1A
1@
1?
1>
1<
1:
19
16
15
11
1,
1+
1*
1(
1'
1&
1%
1$
1HN
1FN
0DN
0BN
0>N
1=N
0<N
08N
15N
11N
0.N
0,N
1%N
1pM
0kM
1jM
1hM
0fM
1dM
1cM
1aM
0`M
1^M
1\M
1[M
0ZM
1YM
0XM
1WM
1VM
0RM
0PM
1MM
1KM
1JM
0FM
1EM
0DM
0BM
0AM
0@M
13M
01M
1/M
0-M
0(M
0&M
1$M
1#M
1~L
0{L
1zL
1]L
1\L
0[L
1ZL
1YL
1WL
0SL
0NL
1LL
0IL
1GL
0CL
0BL
0@L
0?L
1<L
0;L
19L
18L
07L
16L
05L
14L
03L
0/L
1.L
1,L
1+L
0)L
1(L
0PJ
1OJ
0MJ
0HJ
0EJ
0BJ
0>J
0=J
19J
05J
01J
1#J
1~I
0|I
1yI
1jI
1fI
0aI
1]I
1ZI
1YI
0QI
1NI
1LI
0KI
0HI
1>I
1;I
0:I
18I
05I
01I
1dG
1`G
0]G
0\G
0[G
1ZG
1YG
1UG
0SG
0NG
0JG
0GG
1DG
0BG
1@G
1/G
0.G
0,G
0#G
1~F
1}F
0|F
1{F
0wF
1vF
0uF
1tF
0sF
0qF
1pF
1lF
0]F
0ZF
0XF
1VF
1TF
0NF
1LF
1KF
0GF
0EF
0CF
1AF
1=F
0<F
1;F
0:F
09F
18F
06F
05F
1$D
1"D
1}C
1{C
1zC
1xC
1vC
1uC
1sC
1lC
1jC
1iC
1hC
1fC
1dC
1bC
1UC
1TC
1SC
1QC
1NC
1LC
0KC
1FC
1DC
1BC
0AC
1@C
0?C
0=C
1<C
1:C
18C
07C
10C
1.C
0*C
1&C
0$C
1!C
0~B
1xB
0wB
1uB
0sB
0qB
1kB
0cB
0bB
1^B
1]B
1[B
0YB
1WB
1VB
0UB
0TB
1SB
1QB
1PB
0MB
1LB
1HB
1GB
1FB
0DB
0AB
0@B
1?B
0>B
10@
0.@
1-@
1*@
0)@
0(@
1%@
0$@
0~?
0}?
1{?
1x?
1w?
1t?
1q?
0p?
1m?
1b?
0`?
0]?
0\?
1[?
1Y?
1X?
0W?
1V?
0U?
1R?
1P?
0M?
0J?
0I?
0H?
0F?
0E?
1D?
1B?
0A?
0@?
0??
12?
01?
1*?
0)?
1&?
1$?
1"?
0!?
0x>
0h>
0f>
0b>
1a>
0`>
1[>
0Z>
1Y>
1W>
0V>
0R>
1Q>
0P>
0O>
0M>
1J>
0I>
1E>
1D>
1D<
1@<
1=<
0<<
18<
03<
02<
10<
1-<
1,<
0+<
1)<
1&<
0#<
0!<
0z;
0x;
1w;
0v;
0s;
1r;
0q;
1p;
0n;
0l;
0k;
1g;
0d;
1c;
0b;
0a;
0\;
1[;
0Z;
0X;
1W;
1V;
0T;
1S;
0M;
0I;
0H;
0E;
0D;
1B;
0A;
1>;
1<;
09;
06;
02;
1/;
1.;
0&;
1%;
0$;
1#;
1";
1{:
1y:
1x:
0r:
0p:
1o:
1m:
1l:
0k:
1j:
1i:
1d:
0c:
0b:
0a:
0NR
1MR
0LR
1KR
0FR
1CR
0AR
1?R
0>R
0<R
0;R
0:R
17R
05R
14R
1/R
1.R
0-R
1@=
0?=
1>=
0==
0;=
08=
16=
15=
01=
1,=
1*=
0)=
1(=
1'=
0&=
1!=
1~<
0}<
0wR
0uR
0sR
1oR
0nR
1lR
0kR
0iR
1dR
0cR
1bR
0aR
0_R
0^R
1]R
1\R
1[R
1XR
0WR
0VR
0UR
1TR
1PR
14>
10>
0#>
0">
1{=
0y=
1t=
0o=
0vS
0tS
0pS
1iS
0hS
1fS
1eS
0dS
0cS
1aS
0`S
0]S
1[S
0XS
1SS
1RS
13A
12A
01A
0.A
0-A
1,A
1*A
1(A
1'A
0&A
1#A
1"A
0!A
0|@
0y@
0x@
0w@
1t@
1s@
1q@
0p@
1AT
0?T
1>T
1:T
15T
04T
13T
12T
11T
1/T
0.T
1-T
0,T
0+T
0)T
0%T
1#T
0}S
0|S
0{S
1-B
1*B
0(B
1%B
0$B
0~A
0}A
1wA
0CU
0@U
1>U
0=U
0<U
0;U
09U
08U
17U
15U
04U
12U
11U
10U
1-U
0+U
0)U
1(U
0&U
0%U
1$U
0!U
0~T
0|T
1~D
1{D
1yD
1wD
0uD
1tD
1sD
1qD
1pD
0mD
1lD
1hD
0gD
1fD
0eD
0dD
1bD
1`D
1_D
1^D
1hU
1gU
1eU
0aU
0]U
1\U
0[U
0YU
1XU
1VU
1TU
0SU
0QU
1PU
0IU
0HU
1tE
1qE
1lE
1jE
1iE
1^E
0FH
0CH
0AH
0>H
0<H
19H
17H
06H
02H
0/H
1.H
1-H
1*H
1)H
0(H
0$H
0#H
1!H
0~G
1}G
1{G
0yG
1wG
1vH
1tH
0nH
1iH
1fH
0eH
0cH
0`H
1_H
0^H
1]H
0\H
1[H
0ZH
0VH
0:K
17K
15K
04K
13K
11K
10K
0.K
0+K
0)K
0(K
1'K
0&K
1$K
0#K
1zJ
0yJ
1xJ
0vJ
0uJ
0tJ
0qJ
1pJ
0mJ
1lJ
1jJ
1iJ
1hJ
0hK
1bK
1_K
0UK
0QK
1OK
1FK
0EK
0AK
1$W
1#W
0"W
1!W
1~V
1|V
0xV
0vV
0tV
0sV
1rV
0qV
0pV
0nV
1lV
1kV
0iV
1hV
1fV
1eV
0dV
0cV
0aV
0_V
1^V
0]V
0\V
1[V
0ZV
0YV
0XV
0TV
1SV
1QV
1PV
0NV
1MV
1GQ
1FQ
1DQ
1CQ
1AQ
18Q
03Q
11Q
0.Q
0-Q
1,Q
0*Q
1)Q
0(Q
1&Q
0%Q
1$Q
1#Q
0"Q
1!Q
1~P
1}P
1|P
1vP
1tP
1sP
1qP
1pP
1UW
0PW
1OW
1MW
1HW
1GW
1FW
1CW
1>W
1=W
1<W
18W
17W
05W
04W
12W
11W
10W
0+W
1*W
0)W
0(W
0'W
0&W
0%W
1jO
0fO
0`O
1_O
0ZO
0PO
1dP
1cP
1aP
1`P
1^P
1UP
0PP
1NP
0KP
0JP
1IP
0GP
1FP
0EP
1CP
0BP
1AP
1@P
0?P
1>P
1=P
1<P
1;P
15P
13P
12P
10P
1/P
1FX
1EX
0DX
1CX
1BX
1@X
0<X
0:X
08X
16X
05X
04X
11X
10X
1-X
1,X
0'X
1#X
1"X
0!X
1{W
1zW
0xW
1wW
1vW
0tW
0sW
1qW
0oW
0kW
1jW
0iW
0hW
0gW
0fW
0eW
0GQ
0FQ
0DQ
0CQ
0AQ
1;Q
08Q
16Q
01Q
1+Q
1*Q
0)Q
1(Q
1"Q
0!Q
0~P
0}P
0{P
0wP
0vP
0qP
1QD
1ND
1LD
1JD
0HD
1GD
1FD
1DD
1CD
0@D
1?D
1;D
0:D
19D
08D
07D
15D
13D
12D
11D
0=V
0:V
18V
07V
02V
11V
0.V
1,V
1)V
1&V
1%V
1$V
1#V
1!V
0~U
1yU
0xU
0vU
0uU
0tU
1"E
0~D
1}D
0yD
1xD
1uD
0tD
0qD
0pD
1mD
0kD
0aD
0`D
0^D
1a@
1`@
0_@
0\@
0[@
1Z@
1X@
1V@
1U@
0T@
1Q@
1P@
0O@
0L@
0I@
0H@
0G@
1D@
1C@
1A@
0@@
0vT
0tT
0nT
0mT
0hT
0fT
1eT
1bT
1^T
1\T
0ZT
0TT
0ST
0NT
0MT
0LT
03A
0(A
0'A
1&A
1$A
0#A
1y@
0t@
1r<
0q<
1p<
0o<
0m<
0j<
1h<
1g<
0c<
1^<
1\<
0[<
1Z<
1Y<
0X<
1S<
1R<
0Q<
0FS
1ES
1CS
1BS
1@S
0>S
1<S
08S
07S
14S
13S
12S
11S
10S
1.S
0-S
1+S
1*S
0)S
1(S
1'S
0&S
1$S
1#S
0"S
1!S
1{R
0@=
0>=
06=
04=
12=
0/=
0-=
0(=
0'=
0"=
0!=
0~<
0r<
0p<
0h<
0f<
1d<
0a<
0_<
0Z<
0Y<
0T<
0S<
0R<
0l=
1k=
1j=
0g=
1f=
1e=
0d=
0`=
0_=
1^=
0]=
1[=
0Z=
0Y=
0X=
0W=
0R=
0O=
1N=
1M=
1L=
0K=
1H=
1G=
1C=
15>
02>
1->
1,>
0+>
0(>
1'>
1&>
1%>
1$>
1#>
1!>
1}=
1|=
0{=
1z=
1v=
1u=
0t=
0s=
0a@
0V@
0U@
1T@
1R@
0Q@
1I@
0D@
0hA
0fA
1aA
0\A
0[A
0WA
0VA
1UA
0QA
0OA
1NA
1IA
0HA
1GA
0FA
1EA
1DA
1CA
0AA
0?A
0>A
1(B
1'B
0%B
1"B
1!B
0xA
0vA
1pA
0oA
1mA
1SD
0QD
1PD
0LD
1KD
1HD
0GD
0DD
0CD
1@D
0>D
04D
03D
01D
0QE
0NE
1LE
1HE
1EE
0DE
0AE
1>E
08E
07E
13E
02E
11E
1.E
0-E
0*E
0qE
1pE
1mE
1eE
1dE
1cE
1aE
0]E
1[E
1YE
1XE
1VE
0dP
0cP
0aP
0`P
0^P
1XP
0UP
1SP
0NP
1HP
1GP
0FP
1EP
1?P
0>P
0=P
0<P
0:P
06P
05P
00P
1CO
1@O
0>O
1=O
1<O
09O
07O
05O
02O
01O
0-O
1,O
1*O
1(O
1'O
1%O
1#O
1!O
1{N
1zN
0yN
0uN
1tN
1sN
0pN
1oN
0kN
0hN
1gN
0fN
0eN
0dN
0cN
0bN
1$P
1!P
1~O
1sO
1mO
0jO
0hO
0eO
0cO
0]O
1[O
1ZO
1YO
1WO
0VO
1SO
1PO
1MO
1GO
1BO
0AO
1?O
1>O
0<O
06O
13O
11O
0,O
1&O
0%O
0$O
0#O
0{N
0zN
1yN
1xN
1vN
1rN
0qN
0lN
0$P
0!P
0~O
1vO
0sO
1eO
1cO
1]O
0[O
0ZO
0XO
0TO
0ME
0KE
0JE
0FE
0EE
1BE
1AE
0>E
1=E
0:E
18E
0.E
1-E
0+E
1yE
1vE
1qE
0mE
0iE
1fE
0dE
0YE
0aA
1VA
0UA
0TA
0RA
1QA
0IA
0DA
0'B
1%B
1#B
0"B
1xA
0j=
1h=
1`=
0^=
1\=
1Y=
1W=
1R=
1Q=
0L=
1K=
1J=
05>
0->
0&>
0$>
0}=
0|=
0v=
0u=
#54000
b111100111110001100000001 d
b110110101111100110100001101 e
0"
1)Y
0(Y
1'Y
1&Y
0%Y
1!Y
0~X
1}X
1|X
0{X
1xX
0rX
1qX
1pX
0oX
1nX
1mX
0lX
0hX
1u!
0t!
1s!
1r!
0q!
1m!
0l!
1k!
1j!
0i!
1f!
0`!
1_!
1^!
0]!
1\!
1[!
0Z!
0V!
0eX
0bX
0aX
1_X
1^X
0]X
1ZX
1YX
1WX
1SX
1RX
0NX
0KX
0JX
0HX
1G!
0F!
1E!
0C!
0?!
1=!
0<!
1;!
0:!
19!
08!
17!
04!
01!
00!
1/!
0.!
0,!
0+!
0)!
1'!
0%!
0#!
1~
0}
0|
1{
0x
0w
0q
0o
0n
0m
0l
0h
0T!
1r(
0q(
1p(
1o(
0n(
1j(
0i(
1h(
1g(
0f(
1c(
0](
1\(
1[(
0Z(
1Y(
1X(
0W(
0S(
05"
02"
01"
1/"
1."
0-"
1*"
1)"
1'"
1#"
1""
0|!
0y!
0x!
0v!
b0 yQ
b0 vQ
b0 pQ
b0 mQ
b1 jQ
b0 dQ
b1 ^Q
b0 aQ
b1 XQ
b0 RQ
1MQ
1PQ
1VQ
0YQ
1\Q
0_Q
1hQ
0kQ
1tQ
b110110101111100110100001101 KQ
b0 NQ
b0 QQ
b0 TQ
b111111001001010000011001011110010 WQ
b110110101111100110100001101 ZQ
b111110010010100000110010111100101 ]Q
b0 `Q
b0 cQ
b110110101111100110100001101 fQ
b111111001001010000011001011110010 iQ
b0 lQ
b110110101111100110100001101 oQ
b0 rQ
b0 uQ
b0 xQ
1%)
1$)
1")
0!)
1~(
0}(
1z(
0y(
1v(
0q'
0o'
0n'
0l'
0k'
0j'
0i'
0g'
0f'
0d'
0b'
0^'
0['
0Z'
0X'
0W'
0U'
0T'
0S'
0P'
0N'
0M'
0K'
0J'
0I'
0H'
0F'
0E'
0C'
0A'
0='
0:'
09'
07'
06'
04'
03'
02'
0.'
0+'
0&'
0#'
0!'
0}&
0|&
0{&
0y&
0x&
0u&
0r&
0n&
0m&
0g&
0f&
0e&
0_&
1^&
1\&
1[&
1Z&
0Y&
1X&
0P&
0O&
0N&
0K&
0I&
0H&
0F&
0E&
0D&
0C&
0A&
0@&
0>&
0<&
08&
05&
04&
02&
01&
0/&
0.&
0-&
1)&
1&&
1%&
1$&
1#&
1!&
1|%
1{%
1u%
1s%
1p%
1m%
1l%
1k%
1j%
1i%
1h%
1g%
0f%
1e%
1d%
0c%
1_%
0^%
1]%
1\%
0[%
1X%
0R%
1Q%
1P%
0O%
1N%
1M%
0L%
0H%
0G%
0F%
0D%
0C%
0A%
0@%
0?%
0>%
0<%
0;%
09%
07%
03%
00%
0/%
0-%
0,%
0*%
0)%
0(%
0%%
0$%
0"%
0!%
0}$
0|$
0{$
0z$
0x$
0w$
0u$
0s$
0o$
0l$
0k$
0i$
0h$
0f$
0e$
0d$
1b$
1`$
1]$
1\$
1[$
1Z$
1X$
1U$
1T$
1N$
1L$
1I$
1F$
1E$
1D$
1C$
1B$
1A$
0@$
1?$
1>$
0=$
19$
08$
17$
16$
05$
12$
0,$
1+$
1*$
0)$
1($
1'$
0&$
0"$
0!$
1}#
1z#
1y#
1x#
1w#
1u#
1r#
1q#
1k#
1i#
1f#
1c#
1b#
1a#
1`#
1_#
1^#
0[#
0X#
0S#
0P#
0N#
0L#
0K#
0J#
0H#
0G#
0D#
0A#
0=#
0<#
0;#
09#
08#
06#
05#
04#
03#
01#
00#
0.#
0,#
0(#
0%#
0$#
0"#
0!#
0}"
0|"
0{"
0x"
0u"
0p"
0m"
0k"
0i"
0h"
0g"
0e"
0d"
0a"
0^"
0Z"
0Y"
1X"
0W"
1V"
1U"
0T"
1P"
0O"
1N"
1M"
0L"
1I"
0C"
1B"
1A"
0@"
1?"
1>"
0="
09"
08"
08(
1<(
0B(
1@(
0D(
1H(
0J(
0L(
0P(
0R(
0m8
0-,
0,,
0*,
0),
0',
0&,
0%,
0$,
0",
0!,
0}+
0{+
0w+
0t+
0s+
0q+
0p+
0n+
0m+
0l+
1y/
0w/
0v/
0t/
0s/
0q/
0p/
0o/
0n/
0l/
0k/
0i/
0g/
0c/
0`/
0_/
0]/
0\/
0Z/
0Y/
0X/
0+2
0)2
0'2
0&2
0$2
0#2
0"2
0!2
0}1
0|1
0z1
0x1
0t1
0q1
0p1
0n1
0m1
0k1
0j1
0i1
1)5
0'5
0%5
0$5
0"5
0!5
0~4
0}4
0{4
0z4
0x4
0v4
0r4
0o4
0n4
0l4
0k4
0i4
0h4
0g4
0O5
0H5
0G5
0F5
0@5
1?5
1=5
1<5
1;5
0:5
195
015
005
0/5
0#8
0!8
0~7
0|7
0{7
0z7
0y7
0w7
0v7
0t7
0r7
0n7
0k7
0j7
0h7
0g7
0e7
0d7
0c7
0I8
0G8
0E8
0D8
0B8
0A8
0@8
0?8
0=8
0<8
0:8
088
048
018
008
0.8
0-8
0+8
0*8
0)8
0u5
0r5
0o5
0j5
0g5
0e5
0c5
0b5
0a5
0_5
0^5
0[5
0X5
0T5
0S5
1R5
1t2
1q2
1p2
1o2
1n2
1l2
1i2
1h2
1b2
1`2
1]2
1Z2
1Y2
1X2
1W2
1V2
1U2
0T2
0Q2
1O2
0N2
1M2
1L2
0K2
1G2
0F2
1E2
1D2
0C2
1@2
0:2
192
182
072
162
152
042
002
0/2
1.2
1Q/
1O/
1L/
1K/
1J/
1I/
1G/
1D/
1C/
1=/
1;/
18/
15/
14/
13/
12/
11/
00/
1-/
1+/
0*/
1)/
1(/
0'/
1#/
0"/
1!/
1~.
0}.
1z.
0t.
1s.
1r.
0q.
1p.
1o.
0n.
0j.
0i.
1h.
1x,
1u,
1t,
1s,
1r,
1p,
1m,
1l,
1f,
1d,
1a,
1^,
1],
1\,
1[,
1Z,
1Y,
0X,
0U,
0Q,
0N,
0I,
0F,
0D,
0B,
0A,
0@,
0>,
0=,
0:,
07,
03,
12,
00*
0-*
0(*
0%*
0#*
0!*
0~)
0})
0{)
0z)
0w)
0t)
0p)
0o)
1n)
1m)
0l)
1k)
1j)
0i)
1e)
0d)
1c)
1b)
0a)
1^)
0X)
1W)
1V)
0U)
1T)
1S)
0R)
0N)
0M)
0L)
0K)
1J)
1A+
0@+
1?+
0=+
0;+
19+
08+
17+
05+
13+
12+
11+
1/+
0.+
1-+
0,+
0)+
1(+
0&+
0$+
0"+
0!+
0W+
0U+
0S+
0Q+
0D+
0C+
1B+
157
007
0-7
0+7
0*7
1)7
0(7
1{6
0z6
1y6
0w6
0t6
0q6
1n6
0m6
1l6
0[7
0Y7
0V7
0T7
0S7
0Q7
0N7
0L7
0F7
0E7
0C7
0B7
0?7
0=7
0<7
087
074
114
004
0.4
1,4
0+4
1*4
1)4
0(4
0'4
0&4
0%4
1"4
1}3
1|3
1{3
0z3
1x3
0w3
0u3
1t3
1s3
1o3
0n3
0]4
0Z4
1X4
0W4
1S4
0R4
1P4
1M4
1L4
0J4
0G4
0F4
1D4
0C4
1A4
0@4
1:4
191
171
061
151
141
131
021
0/1
0-1
1+1
0*1
0(1
1%1
1#1
0"1
1~0
1}0
1|0
1{0
1z0
0y0
1v0
0t0
1]1
0[1
1W1
1U1
0S1
1P1
0M1
0K1
1I1
0G1
0D1
0@1
1>1
0<1
08.
06.
14.
03.
1/.
1,.
0+.
0*.
0&.
0$.
1".
1~-
0}-
1{-
0z-
1w-
0v-
1s-
0r-
0a.
0].
0Z.
0U.
0M.
0J.
0I.
0F.
0C.
1@.
1>.
0#:
0":
0!:
0}9
0z9
0x9
1w9
0r9
0p9
0n9
1m9
0l9
1k9
1i9
0h9
0f9
0d9
1c9
0K:
0I:
0F:
0D:
0C:
0A:
0?:
0>:
0<:
05:
03:
02:
01:
0/:
0-:
0+:
#55800
1"
1T!
b110110101111100110100001101 N:
b100000000000000000000000000000000000 O:
b101011001001010000011001011110010000000 P:
b10100000000000000000000000000000000000 Q:
b1001011100111110010110010110101001110101 R:
b100000000001000001100001010000010000 S:
b101011000100111011100000110110001010000 T:
b10100001001000000011001001000010000000 U:
b1010100001101101011111001101000011010001 V:
b0 W:
b11110101010101010101010101010000000000 X:
b0 Y:
b100111111011011100001010110001110011011010 "F
b100100011010101000010001000100000 #F
b1000000110101000001100100001010100000101001000 $F
b1001000100110010001010100101001101000000000 %F
b11001100010100101001110001110000110010011000 &F
b101011101011010110001110101101101001000000 'F
b100110110001110110001001100110110010010111000100101001 xK
b101010010101001101001000110100000000 yK
b1111100110110001101011110011010000110011110101000000000 zK
b10000000010000100000100101001000100000000000000000 {K
b10100010100111010110010111000111110001101011000101101111011 HQ
b1000001001001000101001101000101000001010000000010000000000000 IQ
b110100001001110100100000101000000010101010000001101 P!
b10001111010110111000110111110001011110110010001010100100011010 Q!
b111011100100101110100000001001101000001101000101100101001 R!
b10010110100111000101001101000011000000101101011100101101111011 S!
b111100111110001100000001 H!
b10110010110000101000010001100101 J!
b110101110010111101100001101 L!
b10000100100001001101011000001001 N!
b110110101111100110100001101 I!
b10001001001101110101001000010010 K!
b1000110110111111001100110001101 M!
b10110001111100000101011001100011 O!
0iY
1hY
1eY
0dY
0`Y
1\Y
0XY
0WY
1VY
1SY
1RY
0QY
1PY
1MY
1GY
1FY
1EY
1DY
0?Y
0=Y
1<Y
1;Y
18Y
06Y
10Y
1,Y
1c
1b
0a
1`
1_
1]
0Y
0W
0V
1S
0R
0M
1L
0J
0I
0G
1D
0C
0A
0@
0>
1=
0:
17
06
05
13
12
1.
0*
1)
0(
0'
0%
0$
0HN
1BN
1?N
05N
01N
1/N
1&N
0%N
0pM
1mM
1kM
0jM
1iM
1gM
1fM
0dM
0aM
0_M
0^M
1]M
0\M
1ZM
0YM
1RM
0QM
1PM
0NM
0MM
0LM
0IM
1HM
0EM
1DM
1BM
1AM
1@M
16M
14M
0.M
1)M
1&M
0%M
0#M
0~L
1}L
0|L
1{L
0zL
1yL
0xL
0tL
0\L
0YL
0WL
0TL
0RL
1OL
1ML
0LL
0HL
0EL
1DL
1CL
1@L
1?L
0>L
0:L
09L
17L
06L
15L
13L
01L
1/L
1UJ
1RJ
1PJ
1MJ
1LJ
1HJ
1FJ
1BJ
1AJ
1?J
1=J
1:J
09J
17J
14J
12J
0#J
0~I
0}I
1|I
0{I
0zI
1xI
0vI
0tI
1rI
1mI
0jI
0gI
1cI
0bI
1aI
0[I
0ZI
1KI
1HI
1CI
0BI
1AI
1?I
0>I
0=I
17I
06I
10I
0/I
1-I
0fG
0dG
0ZG
0YG
0UG
0RG
0PG
0MG
1LG
0FG
1EG
0DG
1CG
1AG
0?G
0=G
0<G
11G
0/G
1-G
1)G
0(G
0%G
1$G
1"G
0}F
1|F
1wF
0vF
0pF
0lF
0^F
1]F
1ZF
0YF
1XF
1WF
0VF
0QF
0OF
1NF
1MF
0LF
0JF
1CF
0AF
1@F
1?F
1<F
1:F
19F
15F
0$D
0"D
0}C
0{C
0zC
0xC
0vC
0uC
0sC
0lC
0jC
0iC
0hC
0fC
0dC
0bC
0UC
0TC
0SC
0QC
0NC
0LC
1KC
0FC
0DC
0BC
1AC
0@C
1?C
1=C
0<C
0:C
08C
17C
00C
0.C
0+C
0)C
0(C
0&C
0#C
0!C
0yB
0xB
0vB
0uB
0rB
0pB
0oB
0kB
1eB
0`B
0]B
0[B
0ZB
1YB
0XB
1MB
0LB
1KB
0IB
0FB
0CB
1@B
0?B
1>B
00@
0-@
1+@
0*@
1&@
0%@
1#@
1~?
1}?
0{?
0x?
0w?
1u?
0t?
1r?
0q?
1k?
0b?
1\?
0[?
0Y?
1W?
0V?
1U?
1T?
0S?
0R?
0Q?
0P?
1M?
1J?
1I?
1H?
0G?
1E?
0D?
0B?
1A?
1@?
1<?
0;?
14?
02?
1.?
1,?
0*?
1'?
0$?
0"?
1~>
0|>
0y>
0u>
1s>
0q>
1h>
1f>
0e>
1d>
1c>
1b>
0a>
0^>
0\>
1Z>
0Y>
0W>
1T>
1R>
0Q>
1O>
1N>
1M>
1L>
1K>
0J>
1G>
0E>
0D<
0@<
0=<
08<
00<
0-<
0,<
0)<
0&<
1#<
1!<
0w;
0u;
1s;
0r;
1n;
1k;
0j;
0i;
0e;
0c;
1a;
1_;
0^;
1\;
0[;
1X;
0W;
1T;
0S;
0B;
0@;
0>;
0<;
0/;
0.;
1-;
1&;
0%;
1$;
0";
0~:
1|:
0{:
1z:
0x:
1v:
1u:
1t:
1r:
0q:
1p:
0o:
0l:
1k:
0i:
0g:
0e:
0d:
1NR
0MR
1LR
0JR
0HR
1FR
0ER
1DR
0BR
1@R
1>R
1=R
1<R
1:R
06R
15R
03R
01R
0/R
0.R
0,R
0+R
1*R
1A=
1?=
19=
18=
17=
13=
11=
1/=
0.=
1-=
0,=
0*=
1(=
1&=
1$=
1!=
0rR
0oR
1mR
1kR
0gR
0fR
0bR
1^R
0]R
0[R
0XR
1VR
1UR
0TR
0SR
0PR
04>
00>
0~=
0z=
0w=
1o=
1vS
1tS
0sS
1rS
1pS
0lS
0kS
0jS
0iS
1hS
0eS
1dS
1bS
0aS
1`S
1\S
1ZS
1YS
1US
1TS
0SS
0RS
0PS
19A
17A
15A
14A
13A
02A
1-A
0,A
1+A
0*A
1(A
1%A
0$A
1#A
0"A
1~@
1}@
1|@
1{@
1z@
0y@
1w@
1v@
1t@
0s@
0q@
1p@
0AT
0>T
0:T
19T
16T
05T
02T
00T
0/T
1.T
0-T
1,T
1+T
1)T
0&T
1%T
0#T
1"T
1~S
1}S
0xS
00B
0-B
1+B
0*B
1&B
1~A
0{A
0wA
1uA
0tA
1rA
1kA
1EU
0BU
19U
05U
13U
1+U
1*U
0$U
1~T
1|T
1'E
0"E
0}D
0{D
0zD
1yD
0xD
0wD
0rD
1qD
0lD
1kD
0iD
0hD
1gD
0fD
0cD
0bD
1`D
0_D
1^D
0hU
0gU
0eU
1aU
1]U
0\U
1[U
1YU
0XU
0VU
0TU
1SU
1QU
0PU
1IU
1HU
0tE
0nE
0jE
0`E
0^E
0ZE
0XE
0VE
0GH
1FH
1CH
0BH
1@H
0?H
0:H
09H
07H
16H
04H
1/H
1,H
1+H
0*H
0)H
0&H
1#H
0}G
0|G
0{G
1zG
1xG
0vG
0tG
0sG
1xH
0vH
1pH
0oH
1nH
0lH
1kH
0jH
0fH
0bH
1`H
1\H
1UH
14K
03K
01K
00K
1/K
0-K
1)K
0'K
1&K
0%K
0$K
0!K
0~J
0}J
0zJ
1yJ
0xJ
0sJ
0rJ
0pJ
1nJ
0jJ
0iJ
1hK
0fK
1eK
1aK
0]K
1\K
1[K
1XK
1WK
1VK
1QK
1MK
1LK
1JK
1BK
0#W
0~V
0|V
1tV
0rV
1mV
0lV
0jV
0fV
0eV
1dV
1bV
1aV
1`V
1]V
1\V
0[V
1ZV
1YV
1XV
0VV
1TV
19Q
06Q
02Q
11Q
1/Q
1.Q
0,Q
1)Q
0(Q
0$Q
1!Q
1}P
1{P
1wP
1vP
0tP
0sP
0UW
1RW
1PW
0OW
1NW
1LW
1IW
0FW
1EW
0DW
0CW
0AW
1?W
0>W
08W
07W
06W
15W
14W
03W
01W
0.W
1-W
0*W
1(W
1'W
1&W
1%W
1dO
1aO
0WO
0SO
1QO
1HO
0GO
1VP
0SP
0OP
1NP
1LP
1KP
0IP
1FP
0EP
0AP
1>P
1<P
1:P
16P
15P
03P
02P
0EX
0BX
0@X
18X
07X
06X
14X
12X
0+X
1*X
1)X
1'X
1$X
0#X
1}W
0|W
0{W
0zW
0wW
0uW
1tW
1sW
0qW
0nW
1mW
0jW
1hW
1gW
1fW
1eW
09Q
17Q
0/Q
0+Q
0)Q
0&Q
1%Q
0!Q
0wP
1XD
0SD
0PD
0ND
0MD
1LD
0KD
0JD
0ED
1DD
0?D
1>D
0<D
0;D
1:D
09D
06D
05D
13D
02D
11D
1?V
0<V
06V
05V
0-V
0+V
1*V
0)V
0'V
0&V
0%V
1"V
0!V
1}U
1xU
1vU
1uU
1tU
0'E
0yD
0uD
0jD
0`D
0^D
1g@
1e@
1c@
1b@
1a@
0`@
1[@
0Z@
1Y@
0X@
1V@
1S@
0R@
1Q@
0P@
1N@
1M@
1L@
1K@
1J@
0I@
1G@
1F@
1D@
0C@
0A@
1@@
1vT
1tT
0sT
1rT
1mT
1lT
0kT
1jT
0bT
0`T
0_T
0^T
1]T
0[T
1YT
1XT
1ST
1QT
0PT
0OT
1NT
0IT
09A
07A
05A
03A
0/A
1.A
0-A
1,A
0+A
0(A
0#A
0z@
0v@
0u@
0t@
1s@
1s<
1q<
1k<
1j<
1i<
1e<
1c<
1a<
0`<
1_<
0^<
0\<
1Z<
1X<
1V<
1S<
1FS
0ES
1DS
0BS
0@S
0?S
1>S
1=S
16S
05S
03S
02S
1/S
0.S
1-S
0*S
1)S
0(S
0'S
1&S
0%S
0$S
0!S
0~R
0{R
0A=
0?=
09=
08=
07=
05=
01=
0/=
0(=
0&=
0$=
0!=
0|<
1{<
0s<
0q<
0k<
0j<
0i<
0g<
0c<
0a<
0Z<
0X<
0V<
0S<
0P<
1O<
1l=
1j=
0i=
0h=
0f=
0e=
1d=
0b=
0a=
1]=
0\=
0W=
1V=
1U=
1S=
0R=
1O=
0M=
1L=
0J=
0G=
0F=
0C=
16>
10>
1/>
1.>
1)>
0%>
1$>
0#>
0!>
1}=
1q=
0g@
0e@
0c@
0a@
0]@
1\@
0[@
1Z@
0Y@
0V@
0Q@
0J@
0F@
0E@
0D@
1C@
1hA
1gA
1fA
1dA
1cA
0bA
1aA
0`A
1_A
1^A
1]A
1\A
1[A
0ZA
1YA
0XA
0VA
1TA
1SA
1OA
0NA
1LA
1IA
0GA
1FA
0EA
1DA
0BA
0;A
13B
0.B
1'B
0%B
0!B
0~A
1}A
1zA
1yA
0xA
1vA
1tA
0rA
0pA
1oA
0XD
0LD
0HD
0=D
03D
01D
1SE
1RE
0PE
1ME
0IE
0HE
1GE
1FE
1EE
1DE
0AE
0=E
0;E
1:E
08E
14E
10E
1/E
1.E
0-E
1*E
0yE
0vE
0sE
0qE
0pE
0kE
1jE
0fE
0eE
1dE
0aE
0\E
0[E
1YE
1WE
0VP
1TP
0LP
0HP
0FP
0CP
1BP
0>P
06P
0BO
0?O
0=O
15O
03O
0/O
1-O
1,O
0*O
0)O
0(O
0&O
1#O
0!O
0~N
1}N
0yN
1wN
0vN
0tN
1pN
0oN
1kN
1jN
0gN
1eN
1dN
1cN
1bN
1oO
0mO
1jO
1iO
1hO
1fO
0cO
0_O
0YO
1XO
1VO
1SO
0PO
0MO
04O
12O
1*O
1&O
1$O
1!O
1~N
1zN
0rN
0jO
0fO
0dO
0aO
0\O
0RE
0FE
0BE
17E
1-E
1+E
0cE
0YE
0WE
0gA
0eA
0cA
0aA
0]A
0\A
0[A
1ZA
0YA
1VA
0QA
1JA
0FA
1EA
0DA
0CA
1-B
0'B
0yA
0tA
1rA
0k=
1i=
1c=
1b=
1a=
1_=
0[=
0Y=
1R=
0P=
0N=
0K=
0H=
1G=
06>
00>
0/>
0.>
0,>
0}=
#57600
b111011001000111111000101110110 d
b11110100011011100110100111101 e
0"
1%Y
1$Y
0vX
1tX
0sX
0qX
1lX
1kX
1q!
1p!
0d!
1b!
0a!
0_!
1Z!
1Y!
0gX
1fX
1eX
1cX
1bX
1aX
0^X
1[X
0SX
0QX
0PX
1OX
1NX
1LX
1KX
1JX
0G!
1F!
1C!
1?!
1>!
0;!
09!
07!
16!
14!
12!
11!
10!
0-!
1+!
1*!
1(!
0$!
0"!
0!!
0{
1z
1y
1x
1w
1r
1m
1l
1k
0T!
1n(
1m(
0a(
1_(
0^(
0\(
1W(
1V(
07"
16"
15"
13"
12"
11"
0."
1+"
0#"
0!"
0~!
1}!
1|!
1z!
1y!
1x!
0tQ
b1 sQ
0qQ
b1 pQ
1YQ
b0 XQ
0SQ
b1 RQ
0MQ
b1 LQ
b111000010111001000110010110000101 KQ
b111101000110111001101001111010 NQ
b111100001011100100011001011000010 QQ
b111101000110111001101001111010 TQ
b11110100011011100110100111101 WQ
b0 ZQ
b111100001011100100011001011000010 ]Q
b11110100011011100110100111101 fQ
b111000010111001000110010110000101 iQ
b11110100011011100110100111101 lQ
b111100001011100100011001011000010 oQ
b111100001011100100011001011000010 rQ
b11110100011011100110100111101 xQ
0v(
0w(
1!)
0#)
0%)
1q'
1o'
1n'
1m'
1l'
1i'
1g'
1f'
1c'
1b'
1a'
1_'
1^'
1Z'
1X'
1W'
1V'
1U'
1.'
1)'
1('
1&'
1#'
1"'
1|&
1y&
1x&
1w&
1u&
1p&
1o&
1n&
1m&
0l&
1k&
0j&
0i&
1f&
1e&
0d&
1c&
0b&
0a&
1`&
1_&
0^&
0]&
0\&
0Z&
1W&
0U&
1T&
0S&
0R&
1O&
1N&
1M&
1L&
1K&
1I&
1H&
1G&
1F&
1C&
1A&
1@&
1=&
1<&
1;&
19&
18&
14&
12&
11&
10&
1/&
1*&
0)&
1(&
0&&
0%&
0$&
1"&
0!&
1~%
0|%
1z%
1v%
0u%
1r%
1q%
0p%
1o%
0m%
0l%
0k%
1c%
1b%
0V%
1T%
0S%
0Q%
1L%
1K%
0b$
1a$
0`$
0]$
0Z$
1Y$
0X$
1V$
0T$
1Q$
1M$
1J$
0I$
0F$
0A$
0?$
0>$
09$
07$
06$
03$
02$
01$
00$
0/$
0-$
0+$
0*$
0($
0'$
1~#
0}#
1|#
1{#
0x#
0w#
1v#
0u#
1t#
1s#
0r#
0q#
1p#
1o#
1n#
1l#
0i#
1g#
0f#
1e#
1d#
0a#
0`#
0_#
0^#
1\#
1Z#
1Y#
1X#
1W#
1T#
1R#
1Q#
1N#
1M#
1L#
1J#
1I#
1E#
1C#
1B#
1A#
1@#
1;#
16#
15#
13#
10#
1/#
1+#
1(#
1'#
1&#
1$#
1}"
1|"
1{"
1z"
1x"
1v"
1u"
1t"
1s"
1p"
1n"
1m"
1j"
1i"
1h"
1f"
1e"
1a"
1_"
1^"
1]"
1\"
0U"
1Q"
0M"
1K"
0I"
0H"
0G"
0D"
1C"
0>"
1:"
19"
18"
14(
18(
0<(
1L(
1N(
1%8
13*
10*
1.*
1-*
1,*
1+*
1(*
1&*
1%*
1"*
1!*
1~)
1|)
1{)
1w)
1u)
1t)
1s)
1r)
1U,
1R,
1P,
1O,
1N,
1M,
1J,
1H,
1G,
1D,
1C,
1B,
1@,
1?,
1;,
19,
18,
17,
16,
0-/
0+/
0)/
0(/
0#/
0!/
0~.
0{.
0z.
0y.
0x.
0w.
0u.
0s.
0r.
0p.
0o.
0Q/
1P/
0O/
0L/
0I/
1H/
0G/
1E/
0C/
1@/
1</
19/
08/
05/
1K2
1J2
0>2
1<2
0;2
092
142
132
1u2
0t2
1s2
0q2
0p2
0o2
1m2
0l2
1k2
0i2
1g2
1c2
0b2
1_2
1^2
0]2
1\2
0Z2
0Y2
0X2
1'5
1%5
1$5
1#5
1"5
1}4
1{4
1z4
1w4
1v4
1u4
1s4
1r4
1n4
1l4
1k4
1j4
1i4
1G8
1E8
1D8
1C8
1B8
1?8
1=8
1<8
198
188
178
158
148
108
1.8
1-8
1,8
1+8
0j)
1f)
0b)
1`)
0^)
0])
0\)
0Y)
1X)
0S)
1O)
1N)
1M)
1L)
1K)
0J)
1,,
1',
1&,
1$,
1!,
1~+
1z+
1w+
1v+
1u+
1s+
1n+
1m+
1l+
1k+
0j+
1y,
0x,
1w,
1v,
0s,
0r,
1q,
0p,
1o,
1n,
0m,
0l,
1k,
1j,
1i,
1g,
0d,
1b,
0a,
1`,
1_,
0\,
0[,
0Z,
0Y,
1X,
0M5
1L5
0K5
0J5
1G5
1F5
0E5
1D5
0C5
0B5
1A5
1@5
0?5
0>5
0=5
0;5
185
065
155
045
035
105
1/5
1.5
1-5
0,5
1u5
1r5
1m5
1l5
1j5
1g5
1f5
1b5
1_5
1^5
1]5
1[5
1V5
1U5
1T5
1S5
0R5
137
017
0.7
1*7
0)7
1(7
0'7
0#7
0~6
0}6
1|6
0y6
0x6
1w6
0u6
1r6
1q6
1m6
0l6
1Y7
1X7
1V7
1S7
1Q7
1P7
1M7
1L7
1K7
1H7
1D7
1C7
1B7
1A7
1?7
1:7
197
014
104
1.4
0-4
0,4
1+4
0)4
1(4
1'4
1%4
0#4
0"4
1~3
0|3
0{3
1y3
0x3
1w3
1u3
0t3
0s3
1r3
1Y4
0X4
1W4
0S4
1Q4
0P4
0M4
1K4
1B4
0A4
1@4
0<4
091
071
031
001
1/1
0+1
1(1
0&1
0%1
1$1
0#1
1!1
0|0
0z0
0w0
0]1
0W1
0U1
0P1
0O1
0I1
19.
18.
16.
15.
13.
12.
01.
00.
0/.
0,.
1*.
0).
0(.
1#.
1!.
0~-
1}-
1|-
1z-
1y-
0w-
0u-
1t-
0s-
1r-
1[.
1Z.
1Y.
1X.
1U.
1T.
1S.
1P.
1O.
1N.
1M.
1L.
1K.
1D.
1C.
1B.
1A.
0@.
0>.
0A+
1<+
1;+
09+
03+
02+
01+
0/+
1.+
0-+
0++
1%+
1$+
1!+
1~*
1}*
1|*
1e+
1^+
1]+
1X+
1W+
1S+
1P+
1O+
1G+
1F+
0B+
1':
1#:
1!:
1~9
1}9
1|9
0y9
0w9
1v9
0s9
1r9
0q9
0o9
1n9
1j9
1h9
0g9
1f9
0e9
1A:
1?:
1;:
19:
17:
1/:
1-:
#59400
1"
1T!
b111100110110100010100000110001101100 N:
b11000000011001000110000110000001 O:
b1010001111110111000000100010001111101100 P:
b11110000001111110011100111100000000 Q:
b1001011000010111001000110010110000110000 R:
b100000000000000000000000000000000000 S:
b101100101010001110001011011001010010000 T:
b10000010101000000110000100000101000000 U:
b110111000110001100110001010100001000101 V:
b1100001011110001001110011010010110000 W:
b11110010111101100010011000011111010001 X:
b101000000010101000101000000000000 Y:
b10100100101110110000001011111100001101 "F
b10100000000000000001001010000000000000000 #F
b100011011010001101000100011000010101 $F
b101010010011000100100010010100101000001000000 %F
b11111111110110110010100000011101000011010001 &F
b1000001010000000000000000000 'F
b100000011010000111000000011111110000100001000010011010 xK
b100000111011000100001010010100110001000000 yK
b1001101100000001010010000000100100100100101101000000000 zK
b100010001011010100101110111001011001001000000000000000 {K
b1111000111010010010001101011111110110010111001100100101100101001 HQ
b100000000101001010000100000001001101000100000010000000000000 IQ
b11100001110111110001000000110110001111010100000011100011110 P!
b110100001001110100100000101000000010101010000001101 Q!
b10001111010110111000110111110001011110110010001010100100011010 R!
b111011100100101110100000001001101000001101000101100101001 S!
b111011001000111111000101110110 H!
b111100111110001100000001 J!
b10110010110000101000010001100101 L!
b110101110010111101100001101 N!
b11110100011011100110100111101 I!
b110110101111100110100001101 K!
b10001001001101110101001000010010 M!
b1000110110111111001100110001101 O!
1iY
0hY
1gY
0eY
0aY
1_Y
0^Y
1]Y
0\Y
1[Y
0ZY
1YY
0VY
0SY
0RY
1QY
0PY
0NY
0MY
0KY
1IY
0GY
0EY
1BY
0AY
0@Y
1?Y
0<Y
0;Y
05Y
03Y
02Y
01Y
00Y
0,Y
0b
0_
0]
0U
0S
1R
0O
0N
0L
1K
1I
1H
0D
0?
0<
1;
1:
14
03
02
10
1/
0.
1-
0)
0&
1HN
0FN
1EN
1AN
0=N
1<N
1;N
18N
17N
16N
11N
1-N
1,N
1*N
1"N
1jM
0iM
0gM
0fM
1eM
0cM
1_M
0]M
1\M
0[M
0ZM
0WM
0VM
0UM
0RM
1QM
0PM
0KM
0JM
0HM
1FM
0BM
0AM
18M
06M
10M
0/M
1.M
0,M
1+M
0*M
0&M
0"M
1~L
1zL
1sL
0]L
1\L
1YL
0XL
1VL
0UL
0PL
0OL
0ML
1LL
0JL
1EL
1BL
1AL
0@L
0?L
0<L
19L
05L
04L
03L
12L
10L
0.L
0,L
0+L
0UJ
0RJ
0PJ
0OJ
0MJ
0LJ
0JJ
0GJ
0BJ
0AJ
1@J
0?J
0=J
0<J
0:J
08J
07J
06J
04J
02J
1%J
0"J
1}I
0yI
0xI
1wI
1uI
1tI
0rI
0qI
0mI
0kI
1jI
0hI
1gI
1dI
1`I
1_I
1^I
1[I
1ZI
1QI
0NI
0LI
1II
0HI
1DI
0CI
0?I
1=I
0;I
1:I
08I
07I
16I
15I
04I
12I
00I
1/I
1+I
1fG
1dG
0cG
1bG
0`G
0^G
1]G
1\G
0VG
1RG
1QG
0OG
1MG
0LG
1JG
1HG
1GG
0EG
0AG
0@G
09G
01G
0-G
0)G
1&G
0"G
1!G
0~F
0|F
0{F
0wF
0tF
1nF
1lF
1^F
0]F
1\F
0ZF
0XF
0WF
1VF
1UF
1QF
1OF
0NF
0MF
0KF
0IF
1HF
1GF
1EF
0BF
1AF
0@F
0?F
1>F
0=F
0<F
0:F
08F
05F
1xC
1vC
1rC
1pC
1nC
1fC
1dC
1YC
1UC
1SC
1RC
1QC
1PC
0MC
0KC
1JC
0GC
1FC
0EC
0CC
1BC
1>C
1<C
0;C
1:C
09C
1.C
1-C
1+C
1(C
1&C
1%C
1"C
1!C
1~B
1{B
1wB
1vB
1uB
1tB
1rB
1mB
1lB
1cB
0aB
0^B
1ZB
0YB
1XB
0WB
0SB
0PB
0OB
1NB
0KB
0JB
1IB
0GB
1DB
1CB
1?B
0>B
1,@
0+@
1*@
0&@
1$@
0#@
0~?
1|?
1s?
0r?
1q?
0m?
0\?
1[?
1Y?
0X?
0W?
1V?
0T?
1S?
1R?
1P?
0N?
0M?
1K?
0I?
0H?
1F?
0E?
1D?
1B?
0A?
0@?
1??
04?
0.?
0,?
0'?
0&?
0~>
0h>
0f>
0b>
0_>
1^>
0Z>
1W>
0U>
0T>
1S>
0R>
1P>
0M>
0K>
0H>
1><
1=<
1<<
1;<
18<
17<
16<
13<
12<
11<
10<
1/<
1.<
1'<
1&<
1%<
1$<
0#<
0!<
1x;
1w;
1u;
1t;
1r;
1q;
0p;
0o;
0n;
0k;
1i;
0h;
0g;
1b;
1`;
0_;
1^;
1];
1[;
1Z;
0X;
0V;
1U;
0T;
1S;
1P;
1I;
1H;
1C;
1B;
1>;
1;;
1:;
12;
11;
0-;
0&;
1!;
1~:
0|:
0v:
0u:
0t:
0r:
1q:
0p:
0n:
1h:
1g:
1d:
1c:
1b:
1a:
0NR
1MR
1IR
1HR
1ER
0>R
0<R
0:R
07R
12R
11R
1/R
1-R
1,R
1+R
0*R
1<=
1;=
19=
17=
16=
03=
00=
1.=
0-=
1'=
1%=
1$=
1!=
1~<
1}<
1|<
0{<
1uR
1tR
1rR
1qR
1oR
1gR
0eR
0dR
1cR
1bR
1aR
1`R
0^R
1]R
0\R
1[R
1ZR
1XR
0VR
1TR
1RR
1PR
1+>
1(>
1&>
1!>
1u=
1s=
1r=
0q=
0o=
0vS
0tS
1qS
0pS
0mS
1lS
1kS
1iS
0hS
1eS
0dS
0bS
1aS
0`S
1^S
1]S
0[S
0YS
0VS
1/A
0)A
1(A
1'A
0&A
0%A
1$A
1#A
1!A
0}@
0|@
1z@
0w@
1u@
0p@
0;T
09T
07T
06T
15T
14T
03T
1/T
0.T
1-T
1*T
0(T
0'T
0%T
0$T
0"T
0~S
0}S
1|S
1{S
1,B
0+B
1*B
0&B
1$B
0#B
1|A
1sA
1qA
0mA
1CU
0AU
1@U
0?U
0>U
1=U
09U
14U
02U
00U
1.U
0(U
0'U
1&U
1$U
1#U
1!U
0~T
1}T
0|T
1%E
1!E
1zD
1yD
1xD
1wD
1vD
0sD
0qD
1pD
1nD
0mD
0kD
1iD
1hD
1dD
1cD
1bD
1`D
1_D
1kU
1gU
1eU
1dU
1cU
1bU
0_U
1^U
0]U
0YU
0WU
1VU
0UU
1PU
1NU
0MU
0KU
1JU
1fE
1GH
0FH
1EH
0CH
0@H
1>H
1<H
0;H
1:H
18H
06H
15H
14H
0/H
0-H
1'H
1&H
1|G
0xG
0wG
0pG
0xH
1vH
0sH
1rH
0pH
0nH
1mH
0kH
0iH
1hH
1aH
0`H
0_H
0]H
0\H
1WH
0UH
1:K
07K
11K
0/K
1.K
1-K
0,K
1*K
1'K
0&K
1%K
1#K
1!K
0|J
1zJ
0wJ
1sJ
1rJ
1qJ
1pJ
1mJ
1jJ
1iJ
0hK
1fK
0eK
0bK
0aK
0_K
1]K
0\K
0[K
0ZK
0XK
0WK
1UK
0TK
0QK
1PK
0LK
0JK
0FK
0BK
0$W
1#W
1~V
0}V
0zV
0yV
0uV
0tV
1sV
1nV
0mV
1jV
1iV
0gV
1fV
0dV
1cV
0aV
1_V
0^V
0ZV
0YV
1WV
1UV
0SV
0QV
0PV
1FQ
1CQ
1@Q
07Q
16Q
04Q
12Q
1/Q
1-Q
1+Q
0*Q
1'Q
0%Q
0#Q
0"Q
0}P
0|P
0{P
1zP
1xP
1wP
0vP
0pP
1OW
0NW
0LW
1JW
0IW
1BW
1AW
1>W
0<W
09W
17W
16W
05W
04W
1+W
0'W
0&W
0%W
0hO
1^O
1ZO
1YO
1NO
1cP
1`P
1]P
0TP
1SP
0QP
1OP
1LP
1JP
1HP
0GP
1DP
0BP
0@P
0?P
0<P
0;P
0:P
19P
17P
16P
05P
0/P
0FX
1EX
1BX
0AX
0>X
0=X
09X
08X
17X
02X
00X
0-X
0,X
0*X
0(X
0'X
0%X
0$X
0"X
0~W
1{W
0vW
0tW
0sW
1rW
1kW
0gW
0fW
0eW
0FQ
0CQ
13Q
02Q
0/Q
0.Q
1,Q
0+Q
1$Q
1#Q
0xP
1VD
1RD
1MD
1LD
1KD
1JD
1ID
0FD
0DD
1CD
1AD
0@D
0>D
1<D
1;D
17D
16D
15D
13D
12D
1=V
0;V
1:V
08V
17V
15V
12V
01V
00V
1.V
1-V
1+V
0*V
1(V
1'V
1%V
0$V
0#V
0"V
1!V
1~U
0{U
0zU
0xU
0%E
0yD
1rD
0pD
0nD
0gD
0_D
1]@
0W@
1V@
1U@
0T@
0S@
1R@
1Q@
1O@
0M@
0L@
1J@
0G@
1E@
0@@
0vT
0tT
1qT
0pT
0mT
0lT
1kT
0jT
1iT
1fT
1cT
1aT
1`T
0\T
1[T
0WT
1TT
0ST
0QT
1OT
0NT
1MT
1LT
04A
0.A
0(A
0'A
0#A
0~@
0z@
1n<
1m<
1k<
1i<
1h<
0e<
0b<
1`<
0_<
1Y<
1W<
1V<
1S<
1R<
1Q<
1P<
0O<
0FS
1ES
1BS
1@S
1?S
0>S
0=S
0<S
06S
01S
00S
1.S
0-S
0+S
1(S
1$S
1"S
1!S
1}R
1{R
0;=
18=
1*=
0$=
1"=
0m<
1j<
1\<
0V<
1T<
0l=
1k=
1h=
0d=
0b=
0a=
0`=
0]=
1\=
1Z=
1X=
0V=
1T=
0S=
0O=
1K=
0I=
1E=
1C=
13>
12>
1.>
1->
0)>
0'>
0$>
1#>
0!>
1~=
1|=
1z=
1y=
1t=
0r=
0b@
0\@
0V@
0U@
0Q@
0N@
0J@
0hA
0fA
1cA
1bA
0_A
0^A
1\A
1[A
1XA
1WA
0VA
0TA
1QA
0OA
1NA
0LA
0JA
0IA
1GA
1FA
1CA
1AA
1?A
1>A
03B
1.B
0-B
0,B
0(B
1'B
1&B
0$B
1#B
1~A
0|A
1yA
0vA
0uA
0rA
0oA
0VD
0LD
1ED
0CD
0AD
0:D
02D
1QE
1PE
0OE
1NE
1KE
1IE
0GE
0CE
1BE
1AE
1@E
1?E
1=E
0<E
0:E
19E
07E
04E
0/E
0.E
0-E
0,E
1sE
1rE
1oE
0lE
1hE
1gE
1bE
1aE
1`E
1[E
1ZE
1YE
1XE
0cP
0`P
1PP
0OP
0LP
0KP
1IP
0HP
1AP
1@P
07P
0CO
1BO
1AO
1?O
0:O
16O
05O
14O
02O
01O
1)O
1(O
0'O
0&O
0$O
0!O
0~N
0}N
0|N
0wN
1vN
1uN
1rN
0pN
1oN
0kN
1hN
0dN
0cN
0bN
0vO
1qO
0oO
1jO
0iO
1gO
1fO
0eO
1dO
1aO
0ZO
0XO
0QO
1DO
0AO
0>O
0.O
0-O
0*O
0)O
1'O
1&O
1}N
1|N
0sN
1nO
0fO
0PE
1FE
0?E
0=E
1;E
14E
1,E
0rE
1kE
0gE
0`E
0XE
0bA
0\A
1VA
1UA
0QA
0NA
1JA
0'B
0&B
0yA
1e=
1b=
0T=
1N=
0L=
02>
1!>
0y=
1w=
#61200
b1110110110101000101011111101101 d
b1000110001011011111011110001100 e
0"
0)Y
0%Y
0$Y
1"Y
1~X
0|X
1{X
1zX
1rX
0pX
0lX
0kX
1iX
0u!
0q!
0p!
1n!
1l!
0j!
1i!
1h!
1`!
0^!
0Z!
0Y!
1W!
1gX
0fX
1dX
0cX
1`X
1^X
1]X
0ZX
0XX
0WX
0VX
1UX
1SX
0RX
1QX
1PX
0OX
1MX
0LX
1IX
0F!
1@!
0?!
0>!
0=!
19!
18!
15!
13!
02!
01!
1.!
1-!
1,!
0*!
0(!
0'!
1&!
1%!
1!!
0~
1|
1{
0z
0y
0v
1u
0s
0r
1q
1n
0m
0l
0k
1h
0T!
0r(
0n(
0m(
1k(
1i(
0g(
1f(
1e(
1](
0[(
0W(
0V(
1T(
17"
06"
14"
03"
10"
1."
1-"
0*"
0("
0'"
0&"
1%"
1#"
0""
1!"
1~!
0}!
1{!
0z!
1w!
0wQ
b1 vQ
1tQ
b0 sQ
0nQ
b1 mQ
1kQ
b0 jQ
1_Q
b0 ^Q
0PQ
b1 OQ
1MQ
b0 LQ
b1000110001011011111011110001100 KQ
b110111001110100100000100001110011 NQ
b110111001110100100000100001110011 QQ
b0 TQ
b0 WQ
b10001100010110111110111100011000 ZQ
b1000110001011011111011110001100 ]Q
b1000110001011011111011110001100 `Q
b1000110001011011111011110001100 fQ
b1000110001011011111011110001100 iQ
b110111001110100100000100001110011 lQ
b110111001110100100000100001110011 oQ
b10001100010110111110111100011000 rQ
b110111001110100100000100001110011 uQ
b10001100010110111110111100011000 xQ
0u(
1v(
0x(
1y(
1}(
0$)
1%)
0q'
0o'
0l'
1h'
1d'
1`'
0_'
1]'
1['
0Z'
0X'
0U'
1R'
1P'
1O'
1L'
1K'
1J'
1E'
1?'
1<'
1:'
19'
18'
15'
14'
13'
11'
10'
0.'
1,'
1+'
0)'
0('
1''
1%'
1$'
0#'
1!'
1~&
1}&
1z&
0x&
0u&
1s&
1r&
0p&
0o&
0m&
1l&
1h&
1g&
0e&
0c&
1a&
0`&
0_&
0W&
1U&
1Q&
1P&
0N&
1J&
0I&
0H&
1E&
0C&
0A&
0=&
0<&
0;&
1:&
09&
08&
17&
15&
13&
02&
01&
1.&
1,&
1+&
0*&
1'&
1!&
1|%
1y%
1x%
1u%
0r%
0q%
1n%
0i%
0h%
0g%
0c%
0b%
1`%
1^%
0\%
1[%
1Z%
1R%
0P%
0L%
0K%
1I%
1#%
1"%
1|$
1{$
1z$
1y$
1w$
1v$
1u$
1t$
1s$
1q$
1p$
1n$
1j$
1i$
1e$
0a$
1`$
1_$
0\$
1Z$
1X$
1T$
1S$
1R$
0Q$
1P$
1O$
0N$
0L$
0J$
1I$
1H$
0E$
0C$
0B$
1>$
1=$
19$
18$
17$
16$
14$
13$
12$
11$
10$
1.$
1-$
1+$
1'$
1&$
1"$
0~#
0|#
0{#
0z#
0y#
0v#
0t#
0s#
0p#
0o#
0n#
0l#
0k#
0g#
0e#
0d#
0c#
0b#
0\#
0Z#
0Y#
0X#
0W#
0T#
0R#
0Q#
0N#
0M#
0L#
0J#
0I#
0E#
0C#
0B#
0A#
0@#
1<#
18#
17#
05#
03#
11#
00#
0/#
0'#
1%#
1!#
1~"
0|"
1y"
0v"
0p"
0m"
0j"
0i"
0f"
1c"
1b"
0_"
1Z"
1Y"
0X"
1U"
1O"
1L"
1I"
1H"
1E"
0B"
0A"
1>"
09"
08"
04(
16(
0@(
0H(
1J(
0N(
1P(
1/,
1-,
1),
1(,
0&,
0$,
1",
0!,
0~+
0v+
1t+
1p+
1o+
0m+
0R,
0P,
0O,
0N,
0M,
0J,
0H,
0G,
0D,
0C,
0B,
0@,
0?,
0;,
09,
08,
07,
06,
0y,
0w,
0v,
0u,
0t,
0q,
0o,
0n,
0k,
0j,
0i,
0g,
0f,
0b,
0`,
0_,
0^,
0],
1(/
1'/
1#/
1"/
1!/
1~.
1|.
1{.
1z.
1y.
1x.
1v.
1u.
1s.
1o.
1n.
1j.
0y/
1u/
1t/
1p/
1o/
1n/
1m/
1k/
1j/
1i/
1h/
1g/
1e/
1d/
1b/
1^/
1]/
1Y/
0O2
0K2
0J2
1H2
1F2
0D2
1C2
1B2
1:2
082
042
032
112
1O5
1M5
1I5
1H5
0F5
0D5
1B5
0A5
0@5
085
165
125
115
0/5
1I8
0G8
0E8
0B8
1>8
1:8
168
058
138
118
008
0.8
0+8
1(8
0m)
1j)
1d)
1a)
1^)
1])
1Z)
0W)
0V)
1S)
0N)
0M)
0L)
0K)
1J)
03*
11*
0.*
0(*
0%*
0"*
0!*
0|)
1y)
1x)
0u)
1p)
1o)
0n)
0P/
1O/
1N/
0K/
1I/
1G/
1C/
1B/
1A/
0@/
1?/
1>/
0=/
0;/
09/
18/
17/
04/
02/
01/
10/
0u2
1r2
1l2
1i2
1f2
1e2
1b2
0_2
0^2
1[2
0V2
0U2
1T2
0)5
1&5
0%5
0$5
1!5
0}4
0{4
0w4
0v4
0u4
1t4
0s4
0r4
1q4
1o4
1m4
0l4
0k4
1h4
1f4
1e4
0d4
0r5
1p5
1o5
0m5
0l5
1k5
1i5
1h5
0g5
1e5
1d5
1c5
1`5
0^5
0[5
1Y5
1X5
0V5
0U5
0S5
1R5
0%8
1#8
1"8
1}7
1|7
1{7
1v7
1p7
1m7
1k7
1j7
1i7
1f7
1e7
1d7
1b7
1a7
0`7
0?+
0>+
0<+
18+
06+
15+
13+
12+
11+
00+
1/+
0.+
1,+
1++
0*+
1)+
0(+
0'+
0%+
1"+
0!+
0e+
1c+
1b+
0W+
0S+
1R+
0P+
0O+
1L+
1K+
0F+
0':
1$:
0#:
0~9
0}9
0|9
1t9
0r9
1p9
1l9
0j9
1g9
0f9
1e9
1d9
0c9
1K:
1F:
1E:
1@:
1::
15:
13:
1.:
0-:
1+:
057
037
127
107
1.7
0*7
1'7
0&7
1%7
1$7
0"7
0{6
1y6
1x6
0w6
1u6
1o6
0m6
1l6
1[7
0X7
0V7
1U7
1T7
0Q7
0P7
1N7
0M7
0L7
0K7
1J7
1G7
1E7
0B7
0?7
1>7
1=7
1<7
0:7
097
034
114
1/4
1,4
0*4
0'4
1&4
0%4
1"4
0!4
1z3
0y3
1x3
1v3
1s3
1p3
0o3
1n3
0Y4
0W4
1R4
1O4
1M4
1I4
1F4
0D4
0B4
0@4
0:4
051
121
111
101
0.1
0(1
1'1
1&1
0$1
1#1
1"1
0!1
0~0
0}0
1|0
1y0
1x0
1w0
1t0
1r0
1[1
1V1
1U1
1T1
1S1
1R1
1Q1
1P1
1O1
1N1
1M1
1L1
1K1
1I1
1H1
1D1
0>1
1;.
09.
06.
02.
0*.
1(.
1%.
0}-
0y-
1w-
1a.
0[.
0Z.
0Y.
0X.
0U.
0T.
0S.
0P.
0O.
0N.
0M.
0L.
0K.
0D.
0C.
0B.
0A.
#63000
1"
1T!
b111010100001011001011101011001000000 N:
b1000110000010000010000110001100 O:
b1010011011100111010010000010000111001001 P:
b100 Q:
b1011111111011000110011010010011110100000 R:
b100011011111111111100001000000 S:
b1011110111101001101000101001101111000000 T:
b10010111010110000000000000 U:
b1011111001101100100100110110000011101000 V:
b1110010111011010001000011100010100 W:
b11101101110111101000111000010001001000 X:
b10011000101010111000111000110000100 Y:
b101010001001001100100101010010011010011110 "F
b1110100101011010010100101100001000000 #F
b1101010111001001000001011110110000000110000 $F
b100000101000000100110010000001000100000000000 %F
b11111000110110100101000011101110010111100101 &F
b111000001101010101100010001000000000000 'F
b10100111001100011010110011001010101000001101 xK
b1000100000100100010000100001010100000000 yK
b1111111111110000011000010101010110011001101100001000000 zK
b1011000011000000100000000100000000000000000 {K
b1001110010100100110101011001100111000100000001010100100011010 HQ
b1000100000100001001001000110010010010011001001000000000000000000 IQ
b10000010010011011001100100011000011111100111101100000010011100 P!
b11100001110111110001000000110110001111010100000011100011110 Q!
b110100001001110100100000101000000010101010000001101 R!
b10001111010110111000110111110001011110110010001010100100011010 S!
b1110110110101000101011111101101 H!
b111011001000111111000101110110 J!
b111100111110001100000001 L!
b10110010110000101000010001100101 N!
b1000110001011011111011110001100 I!
b11110100011011100110100111101 K!
b110110101111100110100001101 M!
b10001001001101110101001000010010 O!
0iY
1hY
1eY
1aY
1`Y
0]Y
0[Y
0YY
1XY
1VY
1TY
1SY
1RY
0OY
1MY
1LY
1JY
0FY
0DY
0CY
0?Y
1>Y
1=Y
1<Y
1;Y
16Y
11Y
10Y
1/Y
0c
1b
1_
0^
0Z
1V
0R
0Q
1P
1M
1L
0K
1J
1G
1A
1@
1?
1>
09
07
16
15
12
00
1*
1&
0HN
1FN
0EN
0BN
0AN
0?N
1=N
0<N
0;N
0:N
08N
07N
15N
04N
01N
10N
0,N
0*N
0&N
0"N
1pM
0mM
1gM
0eM
1dM
1cM
0bM
1`M
1]M
0\M
1[M
1YM
1WM
0TM
1RM
0OM
1KM
1JM
1IM
1HM
1EM
1BM
1AM
08M
16M
03M
12M
00M
0.M
1-M
0+M
0)M
1(M
1!M
0~L
0}L
0{L
0zL
1uL
0sL
1]L
0\L
1[L
0YL
0VL
1TL
1RL
0QL
1PL
1NL
0LL
1KL
1JL
0EL
0CL
1=L
1<L
14L
00L
0/L
0(L
1OJ
1KJ
0HJ
1GJ
1DJ
1BJ
1>J
1=J
17J
16J
15J
1#J
0!J
1~I
1{I
1yI
0wI
1vI
0sI
1rI
1qI
1pI
0lI
1kI
0jI
1iI
0gI
0_I
0^I
0]I
0QI
1LI
0KI
0II
1HI
0FI
0DI
1>I
06I
05I
13I
02I
11I
0/I
0-I
0fG
0dG
1aG
0]G
0\G
1YG
1VG
1UG
1SG
0RG
0MG
0JG
0GG
1EG
1DG
1AG
1?G
1=G
1<G
10G
1+G
1*G
1(G
0&G
1%G
0$G
1#G
0!G
1~F
1|F
1{F
1yF
1wF
1tF
1rF
1qF
1pF
0nF
0lF
0^F
1]F
1ZF
1WF
0VF
0SF
0RF
0OF
1NF
1LF
1JF
0HF
0EF
0AF
1@F
0>F
1=F
0;F
17F
15F
1$D
1}C
1|C
1wC
1qC
1lC
1jC
1eC
0dC
1bC
0YC
1VC
0UC
0RC
0QC
0PC
1HC
0FC
1DC
1@C
0>C
1;C
0:C
19C
18C
07C
10C
0-C
0+C
1*C
1)C
0&C
0%C
1#C
0"C
0!C
0~B
1}B
1zB
1xB
0uB
0rB
1qB
1pB
1oB
0mB
0lB
0eB
0cB
1bB
1`B
1^B
0ZB
1WB
0VB
1UB
1TB
0RB
0MB
1KB
1JB
0IB
1GB
1AB
0?B
1>B
0,@
0*@
1%@
1"@
1~?
1z?
1w?
0u?
0s?
0q?
0k?
0^?
1\?
1Z?
1W?
0U?
0R?
1Q?
0P?
1M?
0L?
1G?
0F?
1E?
1C?
1@?
1=?
0<?
1;?
12?
1-?
1,?
1+?
1*?
1)?
1(?
1'?
1&?
1%?
1$?
1#?
1"?
1~>
1}>
1y>
0s>
0d>
1a>
1`>
1_>
0]>
0W>
1V>
1U>
0S>
1R>
1Q>
0P>
0O>
0N>
1M>
1J>
1I>
1H>
1E>
1C>
1D<
0><
0=<
0<<
0;<
08<
07<
06<
03<
02<
01<
00<
0/<
0.<
0'<
0&<
0%<
0$<
1z;
0x;
0u;
0q;
0i;
1g;
1d;
0^;
0Z;
1X;
0P;
1N;
1M;
0B;
0>;
1=;
0;;
0:;
17;
16;
01;
0$;
0#;
0!;
1{:
0y:
1x:
1v:
1u:
1t:
0s:
1r:
0q:
1o:
1n:
0m:
1l:
0k:
0j:
0h:
1e:
0d:
0MR
0LR
1JR
0IR
0ER
0CR
1BR
0@R
1>R
0=R
1<R
1:R
19R
16R
05R
13R
02R
0/R
1?=
06=
15=
11=
1/=
0.=
1,=
0*=
1)=
0!=
0}<
1wR
0uR
0tR
0rR
0mR
0lR
0kR
0hR
0gR
1dR
0cR
0bR
0`R
1_R
1^R
0[R
1VR
0TR
14>
0+>
0(>
0&>
0#>
0~=
0|=
0rS
1nS
1mS
0kS
1jS
0iS
1hS
1gS
0fS
1bS
0^S
1[S
1WS
1VS
1SS
1RS
1QS
12A
11A
10A
0/A
1(A
1'A
1&A
1#A
1"A
0!A
1|@
0{@
1y@
1x@
1w@
1v@
0u@
1t@
1r@
0=T
1;T
1:T
19T
18T
16T
04T
13T
01T
0/T
1.T
0,T
0+T
0*T
1'T
1&T
1$T
1#T
1"T
1!T
1}S
1zS
1xS
0*B
1%B
1"B
1wA
0sA
0qA
0kA
0EU
0CU
0@U
1?U
1>U
0=U
1<U
1;U
1:U
18U
06U
03U
01U
0.U
0-U
1,U
0+U
0*U
1'U
0&U
1%U
0$U
0#U
1~T
0}T
1|T
1$E
1~D
0zD
0wD
0vD
1uD
0rD
1nD
1jD
0iD
1gD
1fD
0dD
1aD
1_D
1^D
0kU
0gU
0dU
1]U
1ZU
1XU
1WU
0VU
1MU
1LU
0IU
0HU
1vE
1qE
1pE
1^E
0GH
1FH
1CH
1=H
0<H
17H
05H
04H
12H
00H
1/H
0.H
1-H
0,H
1*H
0'H
0&H
0"H
1~G
0|G
1{G
1xG
1vG
1tG
1sG
1wH
0vH
0tH
1qH
0mH
1lH
1jH
0hH
1gH
1eH
1cH
0aH
1`H
1]H
1YH
0WH
1UH
0:K
05K
04K
13K
02K
10K
1/K
1+K
0)K
0'K
0%K
0#K
1"K
0!K
1~J
1}J
0yJ
1xJ
1wJ
1vJ
1uJ
0oJ
0lJ
1lK
0fK
1_K
1^K
1[K
1ZK
0VK
0UK
1TK
1RK
0PK
0OK
1EK
1$W
0#W
1"W
0~V
0wV
1oV
0nV
1lV
0kV
0jV
0hV
1dV
0cV
1aV
0`V
0_V
1ZV
1YV
0XV
0UV
0TV
0MV
1GQ
1EQ
0@Q
1>Q
0;Q
1:Q
18Q
06Q
15Q
14Q
1/Q
0-Q
1+Q
1(Q
1&Q
1%Q
0$Q
1!Q
1|P
0zP
1xP
1pP
1UW
0RW
1LW
0KW
0JW
0GW
1DW
0AW
0?W
0=W
1<W
0;W
0:W
19W
18W
13W
00W
1.W
1*W
1)W
1'W
1&W
1%W
0jO
1hO
0gO
0dO
0aO
1_O
0^O
0]O
0YO
1WO
0VO
0SO
1RO
0NO
0HO
0DO
1dP
1bP
0]P
1[P
0XP
1WP
1UP
0SP
1RP
1QP
1LP
0JP
1HP
1EP
1CP
1BP
0AP
1>P
1;P
09P
17P
1/P
1FX
0EX
1DX
0BX
0;X
07X
04X
13X
12X
10X
1/X
1-X
0)X
1(X
1'X
0&X
1%X
1$X
1!X
0}W
0yW
1xW
1wW
1vW
1sW
0pW
1oW
1nW
1jW
1iW
1gW
1fW
1eW
0GQ
0EQ
1<Q
04Q
03Q
01Q
0/Q
0(Q
0&Q
0%Q
1}P
0|P
0xP
0wP
0pP
1UD
1QD
0MD
0JD
0ID
1HD
0ED
1AD
1=D
0<D
1:D
19D
07D
14D
12D
11D
0?V
0=V
0:V
18V
07V
16V
14V
10V
0-V
0'V
0!V
0~U
0}U
1|U
1{U
0yU
0wU
0vU
0uU
0tU
1"E
0!E
0~D
1|D
0xD
1qD
1kD
0fD
1eD
1dD
0`D
0_D
1`@
1_@
1^@
0]@
1V@
1U@
1T@
1Q@
1P@
0O@
1L@
0K@
1I@
1H@
1G@
1F@
0E@
1D@
1B@
0rT
1nT
1mT
1lT
0kT
0fT
0eT
0cT
0`T
0]T
1ZT
0YT
1WT
0UT
1PT
1NT
1KT
1IT
01A
00A
1-A
1+A
1*A
1)A
0x@
0w@
1q<
0h<
1g<
1c<
1a<
0`<
1^<
0\<
1[<
0S<
0Q<
0ES
0?S
1=S
0;S
09S
16S
12S
10S
0/S
0.S
0,S
1*S
0(S
1'S
0#S
0!S
0?=
0<=
05=
13=
01=
0/=
1&=
0%=
0q<
0n<
0g<
1e<
0c<
0a<
1X<
0W<
0k=
0i=
0e=
0c=
1a=
1`=
0\=
1[=
1Y=
0U=
1S=
0R=
1P=
0N=
1M=
0K=
0G=
16>
10>
0.>
0->
1)>
1#>
0!>
0t=
0_@
0^@
1[@
1Y@
1X@
1W@
0H@
0G@
0dA
0XA
0WA
0VA
1TA
1RA
1QA
1PA
1HA
0FA
0EA
1DA
1@A
1=A
1;A
11B
10B
1/B
0.B
1'B
0#B
1{A
1xA
1uA
1qA
1SD
0RD
0QD
1OD
0KD
1DD
1>D
09D
18D
17D
03D
02D
0SE
0QE
1OE
0NE
0LE
1JE
1HE
1GE
1CE
0BE
0AE
1?E
17E
06E
15E
12E
1/E
1.E
1-E
0*E
1xE
0vE
0sE
0pE
0oE
1nE
0kE
0aE
1`E
0^E
0[E
1VE
0dP
0bP
1YP
0QP
0PP
0NP
0LP
0EP
0CP
0BP
1<P
0;P
07P
06P
0/P
1CO
1AO
0@O
0?O
0;O
19O
08O
06O
15O
04O
13O
1-O
0,O
0(O
1%O
1$O
0"O
1~N
0}N
0|N
1wN
0vN
1tN
1pN
0mN
1lN
1gN
1fN
1dN
1cN
1bN
1"P
0qO
1pO
1oO
1lO
1jO
1bO
1aO
1^O
1XO
0WO
1UO
0RO
1OO
1MO
0BO
1@O
17O
1/O
1.O
1,O
1*O
0#O
1!O
0~N
0xN
0wN
1sN
0rN
1kN
0"P
0oO
0nO
0lO
0jO
0aO
1ZO
0UO
0MO
0ME
1LE
0KE
0IE
0EE
1>E
18E
03E
02E
01E
0-E
0,E
1yE
0xE
1uE
1^E
1]E
1_A
1^A
0[A
1YA
1XA
1WA
0HA
0GA
00B
0/B
1,B
1i=
1f=
0_=
1]=
0[=
0Y=
0P=
1O=
06>
03>
1{=
0z=
#64800
b1111100111111011110100111111001 d
b11100011001101110010010011000110 e
0"
1(Y
0&Y
1#Y
0!Y
0~X
0{X
0yX
0xX
1vX
0tX
1sX
1oX
0mX
1jX
1hX
1t!
0r!
1o!
0m!
0l!
0i!
0g!
0f!
1d!
0b!
1a!
1]!
0[!
1X!
1V!
0eX
1cX
0^X
0]X
1\X
0[X
1ZX
1XX
1WX
1TX
1RX
0NX
1LX
1F!
0D!
1>!
1<!
1;!
1:!
06!
05!
03!
11!
0/!
0.!
0-!
0,!
1*!
1)!
0&!
0%!
0!!
1}
0|
0{
1z
0w
0u
1p
1o
1m
1i
1g
1f
0T!
1q(
0o(
1l(
0j(
0i(
0f(
0d(
0c(
1a(
0_(
1^(
1Z(
0X(
1U(
1S(
05"
13"
0."
0-"
1,"
0+"
1*"
1("
1'"
1$"
1""
0|!
1z!
b0 vQ
b0 pQ
b1 sQ
b0 mQ
b1 gQ
b1 ^Q
b1 [Q
b0 RQ
0MQ
1PQ
1SQ
0YQ
0eQ
1nQ
1wQ
0zQ
b111100011001101110010010011000110 KQ
b111001100100011011011001110011 NQ
b0 QQ
b111000110011011100100100110001100 WQ
b111001100100011011011001110011 ZQ
b11100110010001101101100111001 ]Q
b0 `Q
b111000110011011100100100110001100 cQ
b11100110010001101101100111001 fQ
b0 iQ
b0 lQ
b111100011001101110010010011000110 oQ
b11100110010001101101100111001 rQ
b0 uQ
b111000110011011100100100110001100 xQ
0%)
1$)
1#)
0!)
0{(
1x(
1u(
0t(
1o'
0m'
1j'
0h'
0g'
0d'
0b'
0a'
1_'
0]'
1\'
1X'
0V'
1S'
1Q'
0P'
0O'
0L'
0K'
0J'
0E'
0?'
0<'
0:'
09'
08'
05'
04'
03'
01'
00'
1/'
1*'
0%'
1#'
0"'
0}&
0|&
0y&
1v&
1q&
0n&
0l&
1j&
0h&
0g&
1e&
1b&
0a&
1_&
1\&
1Z&
1W&
0V&
0U&
1S&
0Q&
0P&
1N&
0K&
0J&
0G&
0F&
0E&
0@&
0:&
07&
05&
04&
03&
00&
0/&
0.&
0,&
0+&
0(&
0'&
0#&
0"&
0!&
0~%
0|%
0{%
0z%
0y%
0x%
0v%
0u%
0s%
0o%
0n%
0j%
1g%
0e%
1c%
1b%
0`%
0]%
1\%
0Z%
0W%
0U%
0R%
1Q%
1P%
0N%
1L%
1K%
0I%
1D%
1C%
1?%
1>%
1;%
18%
15%
14%
13%
11%
10%
1-%
1,%
1(%
1'%
1&%
0#%
0"%
0|$
0{$
0z$
0y$
0w$
0v$
0u$
0t$
0s$
0q$
0p$
0n$
0j$
0i$
0e$
1b$
0`$
1^$
1]$
0[$
0X$
1W$
0U$
0R$
0P$
0M$
1L$
1K$
0I$
1G$
1F$
0D$
1A$
1@$
0>$
1<$
1;$
09$
06$
15$
03$
00$
0.$
0+$
1*$
1)$
0'$
1%$
1$$
0"$
1|#
1{#
1w#
1v#
1s#
1p#
1m#
1l#
1k#
1i#
1h#
1e#
1d#
1`#
1_#
1^#
0<#
0;#
08#
07#
06#
01#
0+#
0(#
0&#
0%#
0$#
0!#
0~"
0}"
0{"
0z"
1p"
1o"
0n"
1m"
1l"
1j"
1i"
0h"
0c"
0Z"
0Y"
1W"
0U"
1R"
0P"
0O"
0L"
0J"
0I"
1G"
0E"
1D"
1@"
0>"
1;"
19"
18"
08(
1>(
1@(
1F(
0J(
1N(
0L(
0P(
0U,
1+/
1*/
0(/
1&/
1%/
0#/
0~.
1}.
0{.
0x.
0v.
0s.
1r.
1q.
0o.
1m.
1l.
0j.
1S/
1Q/
0O/
1M/
1L/
0J/
0G/
1F/
0D/
0A/
0?/
0</
1;/
1:/
08/
16/
15/
03/
1y/
0u/
0t/
0p/
0o/
0n/
0m/
0k/
0j/
0i/
0h/
0g/
0e/
0d/
0b/
0^/
0]/
0Y/
1O2
0M2
1K2
1J2
0H2
0E2
1D2
0B2
0?2
0=2
0:2
192
182
062
142
132
012
1w2
0s2
0r2
0n2
0m2
0l2
0k2
0i2
0h2
0g2
0f2
0e2
0c2
0b2
0`2
0\2
0[2
0W2
0O5
0M5
1K5
0I5
0H5
1F5
1C5
0B5
1@5
1=5
1;5
185
075
065
145
025
015
1/5
0u5
1s5
1n5
0i5
1g5
0f5
0c5
0b5
0_5
1\5
1W5
0T5
0I8
1E8
0C8
1@8
0>8
0=8
0:8
088
078
158
038
128
1.8
0,8
1)8
1'8
0&8
1%8
0#8
0"8
0}7
0|7
0{7
0v7
0p7
0m7
0k7
0j7
0i7
0f7
0e7
0d7
0b7
0a7
1`7
0'5
0&5
0#5
0"5
0!5
0z4
0t4
0q4
0o4
0n4
0m4
0j4
0i4
0h4
0f4
0e4
1d4
1'2
1&2
1"2
1!2
1|1
1y1
1v1
1u1
1t1
1r1
1q1
1n1
1m1
1i1
1h1
1g1
0f1
1w,
1v,
1r,
1q,
1n,
1k,
1h,
1g,
1f,
1d,
1c,
1`,
1_,
1[,
1Z,
1Y,
0X,
0-,
0,,
0),
0(,
0',
0",
0z+
0w+
0u+
0t+
0s+
0p+
0o+
0n+
0l+
0k+
1j+
1(*
1'*
0&*
1%*
1$*
1"*
1!*
0~)
0y)
0p)
0o)
1n)
1l)
0j)
1g)
0e)
0d)
0a)
0_)
0^)
1\)
0Z)
1Y)
1U)
0S)
1P)
1N)
1M)
1L)
1K)
0J)
1@+
1>+
0;+
19+
08+
16+
14+
0/+
1-+
1'+
0$+
0"+
1!+
0b+
1_+
0]+
0X+
1T+
1S+
0R+
0K+
1H+
1F+
1':
0$:
1~9
1z9
1w9
0t9
1q9
0k9
0g9
0d9
0b9
0a9
0`9
0K:
0F:
0E:
0@:
0?:
0::
09:
05:
0.:
1*:
1):
027
0/7
0.7
1,7
0(7
0'7
1&7
0%7
0$7
1#7
0!7
1}6
0|6
1{6
0y6
0x6
0v6
0u6
1s6
0r6
0q6
0p6
0n6
0[7
0Y7
1W7
0U7
0T7
1R7
1O7
0N7
1L7
0J7
1I7
0G7
0E7
0C7
1@7
0>7
0=7
1;7
1:7
134
124
014
0.4
1-4
0,4
0&4
1%4
1#4
0~3
1{3
0z3
1y3
0x3
0u3
1t3
0r3
0q3
1[4
1V4
0Q4
0M4
0K4
0I4
1H4
0F4
1D4
1?4
161
041
131
021
011
0/1
1.1
1+1
1(1
0'1
1~0
0{0
1z0
0y0
0x0
0v0
0u0
0s0
1_1
1]1
0[1
1Z1
1Y1
0V1
0T1
0S1
0Q1
0P1
0N1
0M1
0L1
0K1
0I1
0H1
1G1
0D1
1C1
1B1
08.
05.
04.
12.
1-.
1*.
0(.
1'.
0%.
1$.
0!.
1~-
1}-
0|-
0{-
1y-
0x-
0w-
1v-
1u-
0t-
1s-
0r-
0a.
1>.
#66600
1"
1T!
b111100000101011100011111110100001010 N:
b11100010000001100000000011000100 O:
b101100110011011100100100110001100000001 P:
b10000000000000000000000000000000000000 Q:
b1010100100101010110010110110101001001000 R:
b11000100000001001001000110010100 S:
b1010011011010101001101001001010110110000 T:
b100001000100010010010001000010000 U:
b1001000100000001010001001000001000100000 V:
b111000110010001100100100110001000000 W:
b100110011101100011100110011000001 X:
b1110001000100010001000001000000000000 Y:
b101000000010101010000101001001110001011100 "F
b1010100010000010000010000001000100000 #F
b1011111011000001001001111110111100011000100000 $F
b100010110110110100101000010000100000000 %F
b11010011100011011101001110011011101010010000 &F
b100110011010101010101000100100010001000000 'F
b110101011001101000000110101011000011010011000011110 xK
b100010101001001110100101000011000010000000 yK
b1111011011110111101001101000000011011111010000000000000 zK
b100000001000010100000110111000000000000100000000000 {K
b1111111111100110011100001000010011110010111100010101010000001101 HQ
b10000000010100011001000001001000010000000000000000000 IQ
b1111000111110010001010010000000001110000110010001111101010010110 P!
b10000010010011011001100100011000011111100111101100000010011100 Q!
b11100001110111110001000000110110001111010100000011100011110 R!
b110100001001110100100000101000000010101010000001101 S!
b1111100111111011110100111111001 H!
b1110110110101000101011111101101 J!
b111011001000111111000101110110 L!
b111100111110001100000001 N!
b11100011001101110010010011000110 I!
b1000110001011011111011110001100 K!
b11110100011011100110100111101 M!
b110110101111100110100001101 O!
0hY
1bY
0aY
0`Y
0_Y
1[Y
1ZY
1WY
1UY
0TY
0SY
1PY
1OY
1NY
0LY
0JY
0IY
1HY
1GY
1CY
0BY
1@Y
1?Y
0>Y
0=Y
0:Y
19Y
07Y
06Y
15Y
12Y
01Y
00Y
0/Y
1,Y
1c
0b
1a
0_
0[
1Y
0X
1W
0V
1U
0T
1S
0P
0M
0L
1K
0J
0H
0G
0E
1C
0A
0?
1<
0;
0:
19
06
05
0/
0-
0,
0+
0*
0&
1LN
0FN
1?N
1>N
1;N
1:N
06N
05N
14N
12N
00N
0/N
1%N
0pM
0kM
0jM
1iM
0hM
1fM
1eM
1aM
0_M
0]M
0[M
0YM
1XM
0WM
1VM
1UM
0QM
1PM
1OM
1NM
1MM
0GM
0DM
17M
06M
04M
11M
0-M
1,M
1*M
0(M
1'M
1%M
1#M
0!M
1~L
1{L
1wL
0uL
1sL
0]L
1\L
1YL
1SL
0RL
1ML
0KL
0JL
1HL
0FL
1EL
0DL
1CL
0BL
1@L
0=L
0<L
08L
16L
04L
13L
10L
1.L
1,L
1+L
1UJ
1QJ
0OJ
1MJ
0KJ
1JJ
0GJ
0=J
1<J
1:J
19J
07J
12J
0%J
0#J
1!J
0~I
0}I
0{I
1zI
0yI
1xI
1wI
0uI
1sI
0rI
0qI
1oI
1nI
1hI
1gI
0fI
1eI
0cI
0aI
1_I
1^I
0\I
0ZI
1OI
0LI
1JI
0HI
1EI
1CI
0AI
1@I
1;I
18I
17I
15I
03I
0+I
0bG
1]G
1\G
0YG
1WG
0TG
1RG
1PG
1OG
1NG
0EG
0DG
0CG
1BG
1>G
1;G
19G
11G
00G
1-G
0+G
0*G
0(G
1&G
0%G
0#G
0|F
0{F
0yF
1xF
0wF
0qF
0]F
1XF
0WF
0UF
1SF
1RF
0QF
1OF
0NF
0GF
1EF
0DF
1AF
0@F
1?F
0=F
09F
0$D
0}C
0|C
0wC
0vC
0qC
0pC
0lC
0eC
1aC
1`C
1YC
0VC
1RC
1NC
1KC
0HC
1EC
0?C
0;C
08C
06C
05C
04C
00C
0.C
1,C
0*C
0)C
1'C
1$C
0#C
1!C
0}B
1|B
0zB
0xB
0vB
1sB
0qB
0pB
1nB
1mB
0bB
0_B
0^B
1\B
0XB
0WB
1VB
0UB
0TB
1SB
0QB
1OB
0NB
1MB
0KB
0JB
0HB
0GB
1EB
0DB
0CB
0BB
0@B
1.@
1)@
0$@
0~?
0|?
0z?
1y?
0w?
1u?
1p?
1^?
1]?
0\?
0Y?
1X?
0W?
0Q?
1P?
1N?
0K?
1H?
0G?
1F?
0E?
0B?
1A?
0??
0>?
16?
14?
02?
11?
10?
0-?
0+?
0*?
0(?
0'?
0%?
0$?
0#?
0"?
0~>
0}>
1|>
0y>
1x>
1w>
1e>
0c>
1b>
0a>
0`>
0^>
1]>
1Z>
1W>
0V>
1O>
0L>
1K>
0J>
0I>
0G>
0F>
0D>
0D<
1!<
0w;
0t;
0s;
1q;
1l;
1i;
0g;
1f;
0d;
1c;
0`;
1_;
1^;
0];
0\;
1Z;
0Y;
0X;
1W;
1V;
0U;
1T;
0S;
0M;
1J;
0H;
0C;
1?;
1>;
0=;
06;
13;
11;
1%;
1#;
0~:
1|:
0{:
1y:
1w:
0r:
1p:
1j:
0g:
0e:
1d:
1MR
0KR
0JR
0HR
1GR
0FR
1CR
1AR
1@R
1;R
04R
03R
01R
10R
1/R
1@=
09=
08=
16=
14=
11=
0,=
1+=
0)=
1$=
0"=
1!=
1}<
0|<
0qR
0pR
1nR
1iR
1fR
0dR
1cR
0aR
1`R
0]R
1\R
1[R
0ZR
0YR
1WR
0VR
0UR
1TR
1SR
0RR
0PR
04>
1o=
1pS
0mS
0lS
1kS
0jS
0gS
0bS
0aS
1`S
1_S
0\S
0[S
0ZS
1YS
0VS
0US
0TS
0RS
16A
13A
02A
1/A
1.A
0-A
0*A
0(A
0'A
1}@
1z@
0y@
1w@
0v@
1u@
0t@
1p@
1=T
0;T
08T
06T
12T
10T
1/T
0.T
0-T
1,T
0)T
0&T
0$T
0!T
0|S
0{S
1.B
1)B
0~A
0zA
0wA
1@U
0?U
0;U
19U
08U
07U
04U
10U
0/U
1-U
0,U
1+U
1(U
1#U
0!U
0~T
0$E
1!E
0|D
1xD
1vD
0uD
1tD
1sD
0qD
0nD
1mD
0kD
0jD
0hD
0eD
0dD
0cD
0aD
0^D
1kU
1dU
0cU
0bU
1`U
1\U
0ZU
1VU
1RU
0QU
0MU
1KU
0JU
1HU
0qE
0jE
0dE
0`E
0YE
0FH
0>H
0=H
1<H
1;H
07H
13H
02H
0-H
1)H
1'H
1&H
0#H
1"H
1|G
0{G
0zG
1yG
1uG
1rG
1pG
1xH
0wH
1tH
0rH
0qH
1mH
0jH
0dH
1aH
0`H
1_H
0]H
0YH
0UH
18K
00K
0/K
0-K
0+K
0*K
1(K
1'K
1&K
1%K
1$K
0~J
1|J
0zJ
0xJ
0wJ
0vJ
0uJ
1tJ
0rJ
0pJ
1oJ
1lJ
0jJ
0iJ
0lK
1eK
1cK
1aK
1`K
0_K
0^K
0[K
1XK
1WK
1QK
1PK
1NK
0MK
1IK
0EK
1BK
0$W
1#W
1~V
1zV
1yV
1xV
1tV
1rV
0iV
1gV
0fV
1eV
0dV
1cV
0bV
0aV
1`V
0]V
0\V
1[V
0ZV
0YV
1UV
1SV
1QV
1PV
1FQ
1CQ
1=Q
0<Q
08Q
17Q
05Q
12Q
11Q
00Q
1/Q
1.Q
1-Q
0,Q
1*Q
1)Q
0'Q
0!Q
1~P
0}P
1|P
1{P
1xP
1vP
1tP
1sP
0UW
0PW
1NW
0MW
1KW
1JW
1IW
1FW
0DW
1AW
1@W
0<W
1;W
1:W
09W
08W
07W
06W
14W
0,W
0)W
0(W
0hO
1`O
1]O
1\O
0XO
1TO
1cP
1`P
1ZP
0YP
0UP
1TP
0RP
1OP
1NP
0MP
1LP
1KP
1JP
0IP
1GP
1FP
0DP
0>P
1=P
0<P
1;P
1:P
17P
15P
13P
12P
0FX
1EX
1BX
1>X
1=X
1<X
18X
17X
16X
02X
00X
0/X
1,X
1*X
1)X
0'X
0%X
0$X
1#X
1"X
0!X
1~W
1}W
1zW
1yW
0xW
0vW
1uW
1tW
0sW
0rW
0lW
0iW
0hW
0FQ
0CQ
0>Q
0=Q
07Q
0.Q
1,Q
0*Q
0)Q
1(Q
1!Q
0|P
0UD
1RD
0OD
1KD
1ID
0HD
1GD
1FD
0DD
0AD
1@D
0>D
0=D
0;D
08D
07D
06D
04D
01D
1:V
05V
03V
00V
1)V
0(V
1'V
1&V
0%V
1$V
1"V
1~U
1}U
0{U
1xU
1wU
1vU
1tU
0"E
0!E
1yD
0xD
0tD
1pD
0mD
1kD
1hD
1cD
1aD
1d@
1a@
0`@
1]@
1\@
0[@
0X@
0V@
0U@
1M@
1J@
0I@
1G@
0F@
1E@
0D@
1@@
1pT
0mT
1kT
1eT
1bT
1`T
1^T
1]T
0ZT
1YT
0XT
1VT
0TT
1ST
1RT
0PT
0MT
0LT
03A
10A
0/A
0$A
0#A
0"A
0}@
0z@
0u@
0s@
1r<
0k<
0j<
1h<
1f<
1c<
0^<
1]<
0[<
1V<
0T<
1S<
1Q<
0P<
1ES
0CS
0BS
0@S
1?S
0=S
19S
18S
06S
11S
00S
1.S
1-S
1,S
1+S
0*S
0&S
0$S
1#S
0"S
1!S
1~R
0}R
0{R
0@=
1>=
19=
04=
03=
1.=
0&=
0$=
1#=
0r<
1p<
1k<
0f<
0e<
1`<
0X<
0V<
1U<
1k=
0j=
0i=
0h=
0f=
1e=
0b=
0`=
1_=
1\=
1[=
1W=
1U=
1T=
1R=
0Q=
1P=
1N=
1K=
1J=
1G=
1F=
0E=
0C=
17>
00>
1->
1+>
0)>
0#>
1|=
0{=
0w=
0u=
1t=
0s=
0a@
1^@
0]@
0R@
0Q@
0P@
0M@
0J@
0E@
0C@
1dA
1bA
1aA
1`A
0_A
1\A
1[A
0XA
0WA
1VA
0UA
0TA
0RA
0PA
1OA
0MA
1LA
1KA
1IA
1HA
1GA
1BA
0@A
0?A
0>A
01B
0,B
1(B
0'B
1#B
1!B
1|A
0{A
1yA
0xA
1tA
0qA
1oA
0SD
0RD
1LD
0KD
0GD
1CD
0@D
1>D
1;D
16D
14D
0OE
1NE
0LE
0GE
1EE
0DE
0CE
1BE
1AE
0@E
0>E
1=E
1<E
09E
07E
16E
05E
04E
13E
12E
00E
1-E
1,E
0+E
1*E
1xE
0uE
1oE
0nE
1lE
0hE
0bE
1`E
0^E
0]E
0ZE
0VE
0cP
0`P
0[P
0ZP
0TP
0KP
1IP
0GP
0FP
1EP
1>P
0;P
0CO
1BO
0AO
1?O
1>O
1;O
1:O
09O
18O
07O
05O
14O
12O
10O
0/O
1+O
0*O
1(O
0&O
0%O
0!O
1~N
1}N
1|N
1{N
1yN
1xN
0uN
1rN
0pN
1nN
0iN
0fN
0eN
1#P
1yO
1uO
0pO
0kO
1jO
1iO
1fO
1eO
0bO
1aO
0`O
0_O
0^O
0]O
0\O
0ZO
1YO
1XO
0TO
1SO
1GO
1AO
0>O
19O
08O
02O
1)O
0'O
1%O
0$O
1#O
0zN
1wN
0#P
0yO
0iO
1gO
0eO
1\O
0YO
1ME
1LE
0FE
0EE
0AE
0=E
1:E
08E
15E
10E
0.E
0yE
0xE
1rE
1iE
0fE
1dE
1ZE
0aA
0^A
1]A
1RA
0QA
1PA
1MA
0JA
1EA
0CA
1/B
0.B
0#B
0!B
0|A
0tA
1j=
1h=
1c=
1^=
0]=
0X=
0P=
0N=
0M=
07>
0+>
1%>
1x=
#68400
b11100010111101111000010011000101 d
b11010101000100111101001010101010 e
0"
0'Y
1&Y
1$Y
0#Y
1~X
0}X
1{X
0zX
1yX
1xX
0uX
0rX
0nX
1mX
1kX
0jX
0s!
1r!
1p!
0o!
1l!
0k!
1i!
0h!
1g!
1f!
0c!
0`!
0\!
1[!
1Y!
0X!
1eX
0dX
0cX
0bX
0_X
1]X
0\X
0ZX
0YX
1VX
0TX
1NX
0MX
0LX
0KX
1HX
0E!
1A!
0>!
1=!
0<!
0;!
0:!
16!
15!
04!
12!
1.!
1-!
0+!
0*!
0)!
1(!
1'!
1%!
1$!
1"!
1{
1s
1r
0p
0m
1k
0i
0h
0g
0f
0T!
0p(
1o(
1m(
0l(
1i(
0h(
1f(
0e(
1d(
1c(
0`(
0](
0Y(
1X(
1V(
0U(
15"
04"
03"
02"
0/"
1-"
0,"
0*"
0)"
1&"
0$"
1|!
0{!
0z!
0y!
1v!
1zQ
b1 vQ
1qQ
b1 pQ
0tQ
b0 sQ
b1 jQ
1eQ
0hQ
b0 gQ
b1 aQ
b0 ^Q
0\Q
b0 [Q
b1 UQ
0PQ
b0 OQ
b111010101000100111101001010101010 KQ
b111010101000100111101001010101010 NQ
b101010111011000010110101010101 TQ
b111010101000100111101001010101010 WQ
b111010101000100111101001010101010 ZQ
b0 ]Q
b1010101110110000101101010101011 `Q
b0 cQ
b110101010001001111010010101010100 fQ
b101010111011000010110101010101 iQ
b101010111011000010110101010101 oQ
b111010101000100111101001010101010 rQ
b1010101110110000101101010101011 uQ
b0 xQ
1t(
1w(
0v(
1{(
0z(
0~(
0$)
0o'
0n'
0j'
0i'
0f'
0c'
0`'
0_'
0^'
0\'
0['
0X'
0W'
0S'
0R'
0Q'
1P'
1O'
1M'
1K'
1I'
1G'
1E'
1D'
1B'
1='
1<'
1:'
19'
18'
16'
14'
12'
0/'
1.'
0+'
1('
0''
0$'
1}&
1|&
0z&
1y&
0w&
0v&
1u&
0r&
1o&
1n&
1m&
1l&
0k&
1h&
0e&
1d&
1a&
0\&
0[&
1Y&
0X&
1V&
1U&
0T&
1Q&
0N&
0M&
0L&
1*&
1(&
1&&
1$&
1"&
1~%
1}%
1{%
1v%
1u%
1s%
1r%
1q%
1o%
1m%
1k%
0g%
1e%
0d%
0b%
1a%
0^%
1]%
0\%
0[%
1Z%
0Y%
1W%
1V%
1U%
0T%
1R%
0Q%
0P%
1N%
0M%
0K%
1J%
1H%
1G%
0D%
0C%
0?%
0>%
0;%
08%
05%
04%
03%
01%
00%
0-%
0,%
0(%
0'%
0&%
1%%
1$%
1"%
1~$
1|$
1z$
1x$
1w$
1u$
1p$
1o$
1m$
1l$
1k$
1i$
1g$
1e$
0b$
0_$
0^$
0]$
0Z$
0Y$
0W$
0V$
0T$
0S$
0O$
0L$
0K$
0H$
0G$
0F$
0A$
1>$
0=$
0;$
1:$
07$
04$
13$
10$
0*$
1'$
0&$
0$$
1#$
1"$
1!$
1}#
0|#
1y#
0v#
1u#
0s#
1r#
1o#
1n#
0l#
0k#
1j#
0i#
0h#
1f#
0e#
1b#
1]#
1[#
1Y#
1W#
1U#
1S#
1R#
1P#
1K#
1J#
1H#
1G#
1F#
1D#
1B#
1@#
0y"
1v"
0u"
0s"
1r"
0o"
0l"
1k"
1h"
0b"
1_"
0^"
0\"
1["
1Z"
1Y"
0V"
1U"
1S"
0R"
1O"
0N"
1L"
0K"
1J"
1I"
0F"
0C"
0?"
1>"
1<"
0;"
06(
1:(
0>(
0@(
1B(
0F(
1H(
0N(
1L(
1P(
1)5
0/,
0k)
1j)
1h)
0g)
1d)
0c)
1a)
0`)
1_)
1^)
0[)
0X)
0T)
1S)
1Q)
0P)
1S,
1Q,
1O,
1M,
1K,
1I,
1H,
1F,
1A,
1@,
1>,
1=,
1<,
1:,
18,
16,
1{,
1x,
0w,
1t,
0q,
1p,
0n,
1m,
1j,
1i,
0g,
0f,
1e,
0d,
0c,
1a,
0`,
1],
0S/
0Q/
0N/
0M/
0L/
0I/
0H/
0F/
0E/
0C/
0B/
0>/
0;/
0:/
07/
06/
05/
0y/
1w/
1v/
1t/
1r/
1p/
1n/
1l/
1k/
1i/
1d/
1c/
1a/
1`/
1_/
1]/
1[/
1Y/
0w2
1u2
1s2
1q2
1o2
1m2
1k2
1j2
1h2
1c2
1b2
1`2
1_2
1^2
1\2
1Z2
1X2
0%8
1#8
1"8
1~7
1|7
1z7
1x7
1v7
1u7
1s7
1n7
1m7
1k7
1j7
1i7
1g7
1e7
1c7
01*
1.*
0-*
0+*
1**
0'*
0$*
1#*
1~)
0x)
1u)
0t)
0r)
1q)
1p)
1o)
0n)
0+/
1(/
0'/
0%/
1$/
0!/
0|.
1{.
1x.
0r.
1o.
0n.
0l.
1k.
1j.
1i.
0h.
0O2
1M2
0L2
0J2
1I2
0F2
1E2
0D2
0C2
1B2
0A2
1?2
1>2
1=2
0<2
1:2
092
082
162
052
032
122
102
1/2
0.2
1+2
0'2
0&2
0"2
0!2
0|1
0y1
0v1
0u1
0t1
0r1
0q1
0n1
0m1
0i1
0h1
0g1
1f1
1u5
0s5
1r5
0o5
1l5
0k5
0h5
1c5
1b5
0`5
1_5
0]5
0\5
1[5
0X5
1U5
1T5
1S5
0R5
1M5
0L5
1I5
0F5
1E5
1B5
0=5
0<5
1:5
095
175
165
055
125
0/5
0.5
0-5
1,5
1I8
0E8
0D8
0@8
0?8
0<8
098
068
058
048
028
018
0.8
0-8
0)8
0(8
0'8
1&8
0':
1$:
1":
0!:
1|9
1y9
1x9
0w9
0v9
0u9
1s9
0n9
0m9
0i9
0h9
0e9
1c9
1b9
1a9
1`9
1K:
0A:
1?:
1=:
0;:
15:
11:
1-:
0+:
0*:
0):
174
034
024
004
0/4
0-4
0+4
0(4
1'4
0%4
1!4
0{3
1z3
0w3
0v3
0t3
0s3
1r3
1q3
0p3
0[4
1Y4
1W4
0V4
1U4
1S4
0R4
1Q4
0O4
1N4
0H4
1F4
0D4
1B4
1@4
0?4
1>4
1<4
141
001
0.1
1*1
0(1
1%1
0"1
0|0
0w0
1v0
0t0
1s0
0_1
0]1
0Y1
1X1
1V1
0U1
0R1
1P1
1E1
0B1
1A1
1?1
0>+
09+
07+
04+
03+
01+
1/+
1.+
0,+
0'+
1"+
0!+
0~*
0}*
0|*
0c+
1b+
1`+
0_+
1\+
1W+
1U+
0S+
0L+
1K+
1I+
0H+
0F+
1E+
1D+
1C+
0;.
15.
14.
11.
10.
1/.
1).
1&.
0$.
0#.
0}-
1|-
1{-
1x-
1w-
1_.
1T.
1M.
1L.
1I.
157
007
1/7
1.7
1-7
1+7
1*7
1)7
1(7
1'7
0&7
1$7
1!7
1~6
0}6
0{6
1z6
1x6
1v6
1u6
1t6
1r6
1q6
1p6
1m6
0l6
1Y7
0W7
0S7
0R7
0O7
1N7
0L7
0I7
0H7
1G7
1F7
0D7
1C7
0A7
0@7
0<7
0;7
0:7
187
#70200
1"
1T!
b10000001010111001001100000000010 N:
b11101010100000000110100001010101000 O:
b101111111101010001101100111111111000000 P:
b10000000000100110000001000000000010000 Q:
b1011001000100010010110011110000001101000 R:
b10101010100000001100000101010000000 S:
b1001100000011001011100010000000000000001 T:
b101010100010000010100101010101000000 U:
b101111111101010001101100111111111000001 V:
b10000000000100110000001000000000010000 W:
b11110000000010001101000011111010101000 X:
b101010101010000010100000000000100 Y:
b110011000100111101001110110101010010110 "F
b10000100010001000000100000001000000000000 #F
b1010001101101110111011011001001111100101110000 $F
b10000010001000100100100110000010000000000 %F
b11101101101101100011100100100000101011100000 &F
b10000010001000010010010010000000000000 'F
b101111101100101110001101110001010100001011100000011100 xK
b100010101010100001100000010001000000 yK
b1001111101011000000011001011111000001001010000100000000 zK
b100000010000101110100110100100110101000000000000000000 {K
b1110011011101100111001110111100101001101111010011000011100011110 HQ
b1000000010001000010001000010000110010000000000100000000000000 IQ
b10011011110001011010010110110000110111001101100010011010010 P!
b1111000111110010001010010000000001110000110010001111101010010110 Q!
b10000010010011011001100100011000011111100111101100000010011100 R!
b11100001110111110001000000110110001111010100000011100011110 S!
b11100010111101111000010011000101 H!
b1111100111111011110100111111001 J!
b1110110110101000101011111101101 L!
b111011001000111111000101110110 N!
b11010101000100111101001010101010 I!
b11100011001101110010010011000110 K!
b1000110001011011111011110001100 M!
b11110100011011100110100111101 O!
1hY
0fY
1`Y
1^Y
1]Y
1\Y
0XY
0WY
0UY
1SY
0QY
0PY
0OY
0NY
1LY
1KY
0HY
0GY
0CY
1AY
0@Y
0?Y
1>Y
0;Y
09Y
14Y
13Y
11Y
1-Y
1+Y
1*Y
0c
1b
1_
1[
1Z
0W
0U
0S
1R
1P
1N
1M
1L
0I
1G
1F
1D
0@
0>
0=
09
18
17
16
15
10
1+
1*
1)
0LN
1EN
1CN
1AN
1@N
0?N
0>N
0;N
18N
17N
11N
10N
1.N
0-N
1)N
0%N
1"N
1nM
0fM
0eM
0cM
0aM
0`M
1^M
1]M
1\M
1[M
1ZM
0VM
1TM
0RM
0PM
0OM
0NM
0MM
1LM
0JM
0HM
1GM
1DM
0BM
0AM
18M
07M
14M
02M
01M
1-M
0*M
0$M
1!M
0~L
1}L
0{L
0wL
0sL
0\L
0TL
0SL
1RL
1QL
0ML
1IL
0HL
0CL
1?L
1=L
1<L
09L
18L
14L
03L
02L
11L
1-L
1*L
1(L
0UJ
0QJ
1NJ
0MJ
1KJ
0JJ
1HJ
0FJ
1EJ
0DJ
0BJ
0>J
0:J
09J
05J
02J
0!J
1~I
1}I
0wI
0vI
0tI
0sI
1rI
0pI
0nI
1lI
1jI
0iI
0hI
0gI
1fI
0dI
1cI
1bI
0^I
1]I
1\I
0[I
1ZI
0OI
1MI
0JI
1GI
1FI
0EI
0>I
0;I
0:I
19I
08I
07I
01I
1/I
1bG
1`G
1^G
0]G
0\G
1[G
1ZG
1YG
0VG
0UG
1TG
0SG
0RG
0OG
1MG
1JG
1IG
0HG
1GG
1FG
1EG
1CG
0AG
1@G
0>G
0=G
0<G
01G
0-G
1*G
0&G
1"G
0~F
1yF
0xF
1uF
0tF
0rF
1qF
0pF
1lF
1]F
0[F
0XF
1WF
1UF
0TF
0RF
1QF
1PF
0OF
1NF
1MF
0JF
1IF
1GF
1FF
1DF
0CF
0?F
1=F
1<F
19F
18F
07F
05F
1$D
0xC
1vC
1tC
0rC
1lC
1hC
1dC
0bC
0aC
0`C
0YC
1VC
1TC
0SC
1PC
1MC
1LC
0KC
0JC
0IC
1GC
0BC
0AC
0=C
0<C
09C
17C
16C
15C
14C
1.C
0,C
0(C
0'C
0$C
1#C
0!C
0|B
0{B
1zB
1yB
0wB
1vB
0tB
0sB
0oB
0nB
0mB
1kB
1eB
0`B
1_B
1^B
1]B
1[B
1ZB
1YB
1XB
1WB
0VB
1TB
1QB
1PB
0OB
0MB
1LB
1JB
1HB
1GB
1FB
1DB
1CB
1BB
1?B
0>B
0.@
1,@
1*@
0)@
1(@
1&@
0%@
1$@
0"@
1!@
0y?
1w?
0u?
1s?
1q?
0p?
1o?
1m?
1b?
0^?
0]?
0[?
0Z?
0X?
0V?
0S?
1R?
0P?
1L?
0H?
1G?
0D?
0C?
0A?
0@?
1??
1>?
0=?
06?
04?
00?
1/?
1-?
0,?
0)?
1'?
1z>
0w>
1v>
1t>
1c>
0_>
0]>
1Y>
0W>
1T>
0Q>
0M>
0H>
1G>
0E>
1D>
1B<
17<
10<
1/<
1,<
0z;
1t;
1s;
1p;
1o;
1n;
1h;
1e;
0c;
0b;
0^;
1];
1\;
1Y;
1X;
0N;
1M;
1K;
0J;
1G;
1B;
1@;
0>;
07;
16;
14;
03;
01;
10;
1/;
1.;
0#;
0|:
0z:
0w:
0v:
0t:
1r:
1q:
0o:
0j:
1e:
0d:
0c:
0b:
0a:
1JR
1HR
0GR
1FR
0AR
0@R
0?R
0>R
1=R
0<R
09R
13R
11R
00R
0/R
0>=
09=
15=
14=
13=
1-=
0'=
0#=
1"=
0!=
1|<
0wR
1rR
1qR
1pR
1mR
1lR
1kR
1gR
1eR
1bR
0\R
0[R
1ZR
1YR
1VR
1UR
1sS
1lS
0kS
1jS
1iS
1gS
1fS
0eS
1dS
1bS
0_S
1[S
0YS
1RS
13A
00A
0.A
0+A
1*A
1%A
1#A
0|@
0w@
1v@
1s@
0r@
0p@
1AT
0=T
09T
18T
16T
05T
14T
03T
11T
00T
1+T
1)T
1&T
1%T
0"T
1!T
1|S
0zS
1*B
0)B
1&B
0"B
0yA
0uA
1qA
1mA
1EU
1?U
1=U
1;U
18U
17U
15U
14U
13U
11U
1.U
1,U
0+U
1&U
1$U
1!U
0|T
1'E
1!E
1}D
1|D
1{D
1zD
0yD
1xD
1wD
0vD
1tD
1qD
0pD
0oD
1mD
1lD
1jD
0hD
0gD
1fD
1dD
0cD
0bD
1_D
0kU
1fU
0eU
1bU
1_U
0]U
0[U
1ZU
1YU
0XU
1TU
0SU
0RU
0OU
0KU
1JU
1IU
1jE
1hE
1\E
1FH
0DH
1@H
1>H
08H
16H
15H
14H
12H
1.H
0*H
0'H
0&H
1%H
1$H
0"H
1}G
0|G
1zG
0xG
1wG
0uG
0tG
0sG
0xH
0tH
1qH
1pH
1nH
0mH
0lH
1iH
0eH
1dH
0cH
0_H
1^H
1]H
0[H
1ZH
1YH
1UH
08K
16K
03K
01K
1*K
1)K
0(K
0%K
0$K
0}J
1{J
1zJ
1wJ
1uJ
0tJ
0sJ
1rJ
0qJ
1pJ
0nJ
0mJ
0kJ
1jJ
1iJ
1gK
1fK
0eK
0aK
0`K
0]K
1[K
0ZK
0WK
1UK
0TK
0RK
0QK
0PK
1OK
0NK
1LK
0IK
1FK
0BK
0#W
1{V
0zV
0yV
0xV
1vV
1uV
0tV
0rV
1pV
1nV
1hV
0gV
0cV
1aV
0`V
1^V
1]V
1\V
1YV
0WV
1VV
1RV
1OV
1MV
1<Q
1;Q
13Q
02Q
0-Q
1)Q
0(Q
1'Q
1&Q
1%Q
0#Q
1"Q
1|P
0{P
1zP
1yP
0xP
0vP
1uP
0tP
0sP
1rP
1pP
1SW
0OW
0KW
0JW
0EW
1DW
0@W
1?W
0>W
0:W
19W
17W
15W
02W
10W
0/W
0-W
1)W
1(W
0'W
0&W
0%W
1cO
1bO
0aO
1RO
1PO
0OO
1KO
0GO
1YP
1XP
1PP
0OP
0JP
1FP
0EP
1DP
1CP
1BP
0@P
1?P
1;P
0:P
19P
18P
07P
05P
14P
03P
02P
11P
1/P
0EX
1?X
0>X
0=X
0<X
1:X
19X
08X
06X
15X
14X
12X
01X
0-X
1+X
1&X
1%X
1$X
0{W
0zW
1xW
0wW
0uW
0tW
1rW
1qW
1pW
0mW
1iW
1hW
0gW
0fW
0eW
0;Q
0:Q
03Q
0,Q
0%Q
1#Q
0!Q
0|P
0zP
0yP
0uP
0pP
1XD
1RD
1PD
1OD
1ND
1MD
0LD
1KD
1JD
0ID
1GD
1DD
0CD
0BD
1@D
1?D
1=D
0;D
0:D
19D
17D
06D
05D
12D
1?V
17V
15V
04V
13V
02V
11V
10V
0/V
0.V
0)V
0'V
1%V
0"V
1!V
0|U
1{U
1yU
0wU
1uU
0'E
0!E
0}D
0{D
0wD
1uD
0qD
0lD
0kD
0dD
0aD
1a@
0^@
0\@
0Y@
1X@
1S@
1Q@
0L@
0G@
1F@
1C@
0B@
0@@
1sT
0pT
0kT
1jT
0iT
1hT
1fT
1cT
0`T
0[T
1ZT
0YT
1XT
1UT
1TT
0RT
1QT
1PT
1MT
0KT
06A
0,A
0*A
0)A
0%A
1|@
1z@
0s@
0p<
0k<
1g<
1f<
1e<
1_<
0Y<
0U<
1T<
0S<
1P<
0DS
1BS
1@S
1=S
0:S
17S
16S
15S
02S
01S
1/S
0+S
1&S
0#S
1"S
19=
04=
03=
01=
1/=
1&=
1$=
1k<
0f<
0e<
0c<
1a<
1X<
1V<
0j=
1f=
1`=
0_=
0^=
0\=
0[=
1X=
0U=
1M=
0K=
1I=
0->
1,>
1+>
1*>
1)>
1(>
0%>
1">
0|=
0x=
1w=
0t=
1s=
0d@
0Z@
0X@
0W@
0S@
1L@
1J@
0C@
1eA
0bA
1aA
1^A
0]A
0[A
0ZA
0YA
1UA
0SA
0RA
1QA
0MA
0KA
1JA
0DA
1@A
1?A
0=A
0/B
1,B
1+B
1)B
0&B
1$B
1uA
1sA
1rA
0qA
0oA
0XD
0RD
0PD
0ND
0JD
1HD
0DD
0?D
0>D
07D
04D
1SE
1RE
0LE
1KE
0JE
0BE
1AE
1>E
0<E
0;E
0:E
17E
06E
14E
03E
02E
00E
0-E
0,E
1+E
1xE
1vE
1uE
1sE
0rE
1qE
1pE
0oE
0iE
1fE
1eE
1bE
0`E
1_E
1^E
1]E
1XE
0XP
0WP
0PP
0IP
0BP
1@P
0>P
0;P
09P
08P
04P
0/P
0BO
1<O
0;O
0:O
09O
15O
03O
12O
11O
1/O
0-O
1*O
1$O
0~N
0|N
0{N
0xN
1vN
0sN
0rN
1pN
0kN
0jN
1fN
1eN
0dN
0cN
0bN
1wO
1vO
0uO
0jO
0cO
1aO
1`O
1]O
1ZO
1YO
0XO
1WO
1VO
1TO
0PO
1OO
1MO
1DO
16O
05O
0.O
1'O
1~N
1|N
1zN
0wN
1uN
0tN
0pN
1kN
0vO
0gO
0`O
0\O
0WO
0MO
0RE
1LE
1JE
0HE
1DE
1BE
0>E
19E
18E
11E
1.E
0xE
0vE
0pE
0eE
0dE
0]E
0ZE
0dA
1ZA
1XA
1WA
1SA
0LA
0JA
1CA
0+B
0)B
0(B
0$B
1{A
1yA
0rA
0c=
1^=
1]=
1[=
1Y=
1P=
1N=
10>
0+>
0*>
0(>
#72000
b1110010101011111111011111100101 d
b10111011110100100111001001110111 e
0"
1)Y
1'Y
0&Y
1%Y
1#Y
0"Y
1zX
0xX
0wX
1qX
1pX
1nX
0mX
1lX
1jX
0iX
1u!
1s!
0r!
1q!
1o!
0n!
1h!
0f!
0e!
1_!
1^!
1\!
0[!
1Z!
1X!
0W!
1bX
1_X
1^X
1[X
1ZX
1YX
1TX
0SX
0QX
1KX
0HX
1G!
1B!
0@!
1?!
1;!
1:!
09!
08!
05!
14!
02!
01!
00!
1/!
0.!
1,!
1)!
0(!
0'!
0%!
0$!
1#!
0"!
1!!
1~
0{
1y
0x
1w
1v
0t
0r
1p
0n
1m
0k
1h
1g
1f
0T!
1r(
1p(
0o(
1n(
1l(
0k(
1e(
0c(
0b(
1\(
1[(
1Y(
0X(
1W(
1U(
0T(
12"
1/"
1."
1+"
1*"
1)"
1$"
0#"
0!"
1y!
0v!
0zQ
b1 mQ
1hQ
b0 aQ
b1 ^Q
1YQ
b1 RQ
b0 UQ
b110111011110100100111001001110111 KQ
b110111011110100100111001001110111 NQ
b10001000010110110001101100010001 QQ
b0 TQ
b0 WQ
b101110111101001001110010011101110 ZQ
b1000100001011011000110110001000 ]Q
b0 `Q
b0 fQ
b1000100001011011000110110001000 iQ
b1000100001011011000110110001000 lQ
b1000100001011011000110110001000 oQ
b110111011110100100111001001110111 rQ
b1000100001011011000110110001000 uQ
b101110111101001001110010011101110 xQ
0t(
1z(
1!)
1p'
1o'
1n'
1l'
1k'
1j'
1g'
1d'
1c'
1b'
1_'
1\'
1Z'
1Y'
1X'
1W'
1U'
1T'
1S'
1Q'
0P'
0O'
0K'
1H'
0G'
1F'
0D'
0B'
1A'
1@'
1>'
0<'
1;'
0:'
09'
08'
04'
1/'
1-'
0,'
1+'
1)'
0('
1"'
0~&
0}&
1w&
1v&
1t&
0s&
1r&
1p&
0o&
0l&
0j&
1i&
0h&
0f&
1e&
0_&
1]&
1\&
0V&
0U&
0S&
1R&
0Q&
0O&
1N&
1H&
1D&
1C&
1A&
1@&
1<&
1;&
19&
18&
16&
11&
1-&
0*&
0(&
1'&
0&&
0$&
1#&
0{%
1y%
1x%
0r%
0q%
0o%
1n%
0m%
0k%
1j%
0e%
0c%
0a%
0_%
0]%
0Z%
0X%
0W%
0V%
0U%
0R%
0N%
0L%
0J%
0H%
0G%
0%%
0$%
0"%
0~$
0|$
0z$
0x$
0w$
0u$
0p$
0o$
0m$
0l$
0k$
0i$
0g$
0e$
1_$
1[$
1Z$
1X$
1W$
1S$
1R$
1P$
1O$
1M$
1H$
1D$
1?$
1;$
08$
17$
05$
14$
01$
00$
1/$
0-$
1,$
1*$
1($
1$$
0"$
0}#
0{#
0y#
0w#
0u#
0r#
0p#
0o#
0n#
0m#
0j#
0f#
0d#
0b#
0`#
0_#
0^#
0]#
0[#
0Y#
0W#
0U#
0S#
0R#
0P#
0K#
0J#
0H#
0G#
0F#
0D#
0B#
0@#
1<#
18#
14#
13#
11#
10#
1,#
1+#
1)#
1(#
1&#
1!#
1{"
1y"
1w"
0v"
1u"
1s"
0r"
1l"
0j"
0i"
1c"
1b"
1`"
0_"
1^"
1\"
0["
1X"
1V"
0U"
1T"
1R"
0Q"
1K"
0I"
0H"
1B"
1A"
1?"
0>"
1="
1;"
0:"
0:(
18(
1@(
0B(
1J(
0+2
1m)
1k)
0j)
1i)
1g)
0f)
1`)
0^)
0])
1W)
1V)
1T)
0S)
1R)
1P)
0O)
11*
1/*
0.*
1-*
1+*
0**
1$*
0"*
0!*
1y)
1x)
1v)
0u)
1t)
1r)
0q)
1-,
1),
1%,
1$,
1",
1!,
1{+
1z+
1x+
1w+
1u+
1p+
1l+
1U,
0S,
0Q,
0O,
0M,
0K,
0I,
0H,
0F,
0A,
0@,
0>,
0=,
0<,
0:,
08,
06,
1)/
1%/
0"/
1!/
0}.
1|.
0y.
0x.
1w.
0u.
1t.
1r.
1p.
1l.
0j.
1N/
1J/
1I/
1G/
1F/
1B/
1A/
1?/
1>/
1</
17/
13/
1y/
0w/
0v/
0t/
0r/
0p/
0n/
0l/
0k/
0i/
0d/
0c/
0a/
0`/
0_/
0]/
0[/
0Y/
0u2
0s2
1r2
0q2
0o2
1n2
0h2
1f2
1e2
0_2
0^2
0\2
1[2
0Z2
0X2
1W2
1$5
1~4
1}4
1{4
1z4
1v4
1u4
1s4
1r4
1p4
1k4
1g4
1O5
0M5
0K5
1J5
0I5
0G5
1F5
0@5
1>5
1=5
075
065
045
135
025
005
1/5
1s5
1q5
0p5
1o5
1m5
0l5
1f5
0d5
0c5
1]5
1\5
1Z5
0Y5
1X5
1V5
0U5
0#8
0"8
0|7
1y7
0x7
1w7
0u7
0s7
1r7
1q7
1o7
0m7
1l7
0k7
0j7
0i7
0e7
0{,
0x,
0v,
0t,
0r,
0p,
0m,
0k,
0j,
0i,
0h,
0e,
0a,
0_,
0],
0[,
0Z,
0Y,
1X,
0M2
0K2
0I2
0G2
0E2
0B2
0@2
0?2
0>2
0=2
0:2
062
042
022
002
0/2
1.2
1F8
1E8
1D8
1B8
1A8
1@8
1=8
1:8
198
188
158
128
108
1/8
1.8
1-8
1+8
1*8
1)8
1'8
0&8
1%:
0$:
0":
1!:
0|9
0y9
1u9
1r9
0q9
1n9
1m9
1k9
1j9
1i9
1h9
1e9
1d9
0c9
0a9
0`9
0K:
1H:
1D:
1C:
1A:
0=:
1<:
1;:
19:
05:
03:
1+:
1):
137
117
107
0.7
0+7
0*7
0#7
1}6
1|6
1y6
0x6
0u6
0q6
0p6
0o6
0Y7
1V7
1S7
1R7
1Q7
1K7
1J7
1I7
0G7
0C7
1A7
1?7
1;7
1:7
031
111
101
1.1
0,1
0*1
1(1
0%1
0~0
1}0
1|0
1{0
0z0
1x0
1w0
0v0
0s0
1]1
0X1
0V1
1U1
1R1
0P1
0O1
1M1
1J1
1H1
0G1
0E1
0A1
04.
03.
02.
0/.
0*.
1(.
0'.
1%.
1#.
0".
0~-
0{-
0z-
0y-
0w-
0u-
1t-
0s-
1r-
1a.
0_.
0T.
0M.
0L.
0I.
0>.
1A+
1>+
1<+
1:+
19+
18+
14+
11+
10+
0/+
0++
1*+
0)+
1'+
1%+
1#+
0"+
1!+
1c+
0b+
1a+
0`+
1_+
0^+
0\+
0U+
0T+
1O+
1M+
1L+
0K+
1J+
0I+
1H+
0G+
1F+
0E+
074
1.4
1*4
1)4
1&4
0#4
1|3
0y3
1u3
1p3
0Y4
0W4
0U4
0S4
0Q4
0N4
0L4
0F4
0B4
0@4
0>4
0<4
#73800
1"
1T!
b101010100100110111011101110101011 N:
b11010101011010000000100000001010100 O:
b1010101000100001011011000110110001000000 P:
b100 Q:
b1010000110011100010010110100101100101000 R:
b10001000010100100001001000010010000 S:
b1011100100001011011000110110001000000000 T:
b0 U:
b100001110100110111100100111001101110101 V:
b10110001010000100111001001110010000000 W:
b101100111111101011010010110011000100 X:
b1010101010000010101100101011000100000 Y:
b110110011110111001111101101100011010010 "F
b10001000100000000100000010010001000000000 #F
b1000111110101110000011101011110101010110101000 $F
b1000001010001010100000100001010000000000000 %F
b11110011010011011100000101101000001111100001 &F
b1000101100100010101010000101010000000000 'F
b101000110110011100110001010011011111100011101010010110 xK
b100011001100100100101000010110000000000000 yK
b1110100110100101001110001000110110001000000010000000000 zK
b10000010010000010010010000000100110000000000000000 {K
b1111001101100000110011011100111011111100111101010000010011100 HQ
b1000000100010011101001100100011000100000000000000001000000000000 IQ
b1110000101110100110110011101000001001101000010100011010101110011 P!
b10011011110001011010010110110000110111001101100010011010010 Q!
b1111000111110010001010010000000001110000110010001111101010010110 R!
b10000010010011011001100100011000011111100111101100000010011100 S!
b1110010101011111111011111100101 H!
b11100010111101111000010011000101 J!
b1111100111111011110100111111001 L!
b1110110110101000101011111101101 N!
b10111011110100100111001001110111 I!
b11010101000100111101001010101010 K!
b11100011001101110010010011000110 M!
b1000110001011011111011110001100 O!
0gY
1cY
0`Y
1_Y
0^Y
0]Y
0\Y
1XY
1WY
0VY
1TY
1PY
1OY
0MY
0LY
0KY
1JY
1IY
1GY
1FY
1DY
1?Y
17Y
16Y
04Y
01Y
1/Y
0-Y
0,Y
0+Y
0*Y
0b
1\
0[
0Z
0Y
1U
1T
1Q
1O
0N
0M
1J
1I
1H
0F
0D
0C
1B
1A
1=
0<
1:
19
08
07
04
13
01
00
1/
1,
0+
0*
0)
1&
1GN
1FN
0EN
0AN
0@N
0=N
1;N
0:N
07N
15N
04N
02N
01N
00N
1/N
0.N
1,N
0)N
1&N
0"N
0nM
1lM
0iM
0gM
1`M
1_M
0^M
0[M
0ZM
0UM
1SM
1RM
1OM
1MM
0LM
0KM
1JM
0IM
1HM
0FM
0EM
0CM
1BM
1AM
08M
04M
11M
10M
1.M
0-M
0,M
1)M
0%M
1$M
0#M
0}L
1|L
1{L
0yL
1xL
1wL
1sL
1\L
0ZL
1VL
1TL
0NL
1LL
1KL
1JL
1HL
1DL
0@L
0=L
0<L
1;L
1:L
08L
15L
04L
12L
00L
1/L
0-L
0,L
0+L
1QJ
1OJ
0NJ
1MJ
0KJ
1FJ
0EJ
1DJ
1BJ
0@J
1>J
0<J
1;J
1:J
18J
06J
14J
1%J
1{I
0xI
1tI
1qI
0lI
0kI
0jI
1iI
1hI
1gI
0fI
1dI
0cI
0bI
1aI
0`I
1^I
0]I
0\I
1[I
0MI
1JI
1HI
0GI
0FI
0@I
1;I
13I
0/I
1-I
1cG
0bG
0`G
1_G
1\G
0[G
0YG
0WG
1VG
1UG
1SG
0PG
1OG
0KG
0JG
0IG
0BG
1AG
1>G
1=G
0;G
1-G
0*G
1)G
1&G
0"G
1}F
0yF
0uF
1tF
0qF
1pF
0\F
1XF
0UF
1RF
0QF
1OF
0NF
1KF
1JF
0GF
1BF
1@F
1?F
0=F
1;F
0$D
1!D
1{C
1zC
1xC
0tC
1sC
1rC
1pC
0lC
0jC
1bC
1`C
1WC
0VC
0TC
1SC
0PC
0MC
1IC
1FC
0EC
1BC
1AC
1?C
1>C
1=C
1<C
19C
18C
07C
05C
04C
0.C
1+C
1(C
1'C
1&C
1~B
1}B
1|B
0zB
0vB
1tB
1rB
1nB
1mB
1cB
1aB
1`B
0^B
0[B
0ZB
0SB
1OB
1NB
1KB
0JB
0GB
0CB
0BB
0AB
0,@
0*@
0(@
0&@
0$@
0!@
0}?
0w?
0s?
0q?
0o?
0m?
0b?
1Y?
1U?
1T?
1Q?
0N?
1I?
0F?
1B?
1=?
14?
0/?
0-?
1,?
1)?
0'?
0&?
1$?
1!?
1}>
0|>
0z>
0v>
0b>
1`>
1_>
1]>
0[>
0Y>
1W>
0T>
0O>
1N>
1M>
1L>
0K>
1I>
1H>
0G>
0D>
1D<
0B<
07<
00<
0/<
0,<
0!<
0s;
0r;
0q;
0n;
0i;
1g;
0f;
1d;
1b;
0a;
0_;
0\;
0[;
0Z;
0X;
0V;
1U;
0T;
1S;
1N;
0M;
1L;
0K;
1J;
0I;
0G;
0@;
0?;
1:;
18;
17;
06;
15;
04;
13;
02;
11;
00;
1&;
1#;
1!;
1}:
1|:
1{:
1w:
1t:
1s:
0r:
0n:
1m:
0l:
1j:
1h:
1f:
0e:
1d:
1NR
0JR
0HR
1ER
0DR
1AR
1>R
08R
06R
15R
03R
01R
0-R
1A=
1>=
1<=
1:=
18=
07=
06=
14=
11=
0/=
0.=
0+=
1*=
1)=
1'=
0&=
1%=
0$=
1#=
0"=
1!=
0~<
0}<
1tR
0rR
0pR
0oR
0nR
0kR
0gR
0fR
1dR
0cR
1aR
0`R
0^R
0YR
0XR
0WR
0UR
0SR
1RR
1PR
14>
0o=
0qS
0pS
0nS
1mS
0lS
1kS
0jS
0gS
0fS
1eS
0dS
1cS
0bS
1aS
1^S
0]S
1ZS
0WS
1VS
0RS
03A
10A
1.A
1*A
1(A
1%A
1}@
1{@
0z@
1x@
1w@
0v@
0AT
0:T
06T
13T
02T
10T
0/T
1(T
0'T
0%T
0#T
0}S
1{S
1zS
0,B
0*B
0}A
0sA
0mA
1CU
1AU
0>U
0=U
0;U
09U
08U
03U
12U
01U
00U
1/U
1+U
0(U
0'U
0&U
0#U
1%E
1#E
1}D
0|D
0zD
1yD
0sD
1oD
1lD
1kD
0jD
1hD
1gD
1eD
1dD
1cD
1bD
1iU
0fU
0bU
0aU
0`U
0_U
0^U
1[U
0ZU
0YU
0WU
0VU
0TU
1SU
1RU
1QU
1OU
0NU
1KU
0JU
0IU
0HU
0GU
1oE
1nE
0hE
1gE
0^E
0EH
1AH
0>H
1=H
0<H
17H
06H
05H
03H
0.H
1,H
1'H
0yG
1xG
1uG
1tG
0rG
1sH
0qH
1oH
0nH
1mH
1lH
1jH
0iH
0gH
1fH
1eH
1_H
0^H
0ZH
06K
15K
13K
11K
10K
1/K
1-K
0)K
1(K
0'K
1#K
1}J
1xJ
0uJ
0pJ
0oJ
1nJ
0lJ
0gK
0fK
1]K
0UK
1RK
0OK
1NK
1MK
0LK
1JK
1HK
0FK
1DK
1#W
0!W
1yV
1wV
1tV
1mV
0lV
1iV
0hV
1gV
1fV
0eV
1_V
0^V
0\V
1ZV
0YV
1XV
1WV
0UV
1TV
0RV
0QV
0PV
1FQ
1>Q
16Q
14Q
12Q
01Q
1.Q
0'Q
0&Q
1%Q
1$Q
0#Q
0"Q
1}P
1zP
1yP
1xP
1wP
1uP
1sP
0rP
1pP
0SW
1QW
0NW
0LW
1JW
0IW
0HW
1EW
0?W
1>W
1=W
05W
03W
00W
0.W
1-W
1,W
0+W
0*W
0)W
0(W
1'W
1&W
1%W
0YO
0VO
0TO
0SO
0RO
0KO
0DO
1cP
1[P
1SP
1QP
1OP
0NP
1KP
0DP
0CP
1BP
1AP
0@P
0?P
1<P
19P
18P
17P
16P
14P
12P
01P
1/P
1EX
0CX
1=X
1;X
18X
05X
03X
11X
0.X
1-X
0)X
1'X
0#X
0"X
1!X
0}W
1|W
1{W
1zW
0yW
1wW
1vW
1uW
1tW
0rW
0pW
0nW
1mW
1lW
0kW
0jW
0iW
0hW
1gW
1fW
1eW
0FQ
0>Q
0<Q
02Q
11Q
0.Q
1,Q
0+Q
1!Q
0}P
0xP
0wP
0uP
0sP
1VD
1TD
1PD
0OD
0MD
1LD
0FD
1BD
1?D
1>D
0=D
1;D
1:D
18D
17D
16D
15D
1=V
1;V
08V
05V
14V
03V
12V
00V
1/V
1.V
0+V
1*V
1(V
1'V
0$V
0}U
1zU
1wU
0vU
0uU
0tU
0sU
0%E
0#E
1rD
1qD
1pD
0kD
0gD
0cD
0a@
1^@
1\@
1X@
1V@
1S@
1M@
1K@
0J@
1H@
1G@
0F@
0qT
0nT
1mT
0lT
1kT
0jT
1iT
1gT
0fT
0dT
0cT
1_T
0]T
0ZT
0TT
0NT
1LT
1KT
14A
11A
00A
0.A
0*A
1)A
0(A
0%A
0w@
1s<
1p<
1n<
1l<
1j<
0i<
0h<
1f<
1c<
0a<
0`<
0]<
1\<
1[<
1Y<
0X<
1W<
0V<
1U<
0T<
1S<
0R<
0Q<
1FS
0BS
1AS
0@S
0?S
1;S
09S
08S
06S
04S
13S
11S
0)S
0&S
1$S
0"S
0~R
1}R
1{R
0A=
08=
0)=
0s<
0j<
0[<
1l=
0k=
1g=
0e=
1d=
1b=
0`=
1_=
1\=
0[=
0Z=
0X=
0W=
1U=
0T=
0S=
1Q=
0P=
0N=
0M=
1K=
0I=
1H=
0F=
1E=
1C=
18>
04>
0,>
0)>
1(>
1$>
0">
1!>
1~=
1x=
0w=
0s=
1b@
1_@
0^@
0\@
0X@
1W@
0V@
0S@
0G@
0cA
0aA
0`A
1_A
1]A
1[A
1YA
0UA
0SA
0QA
0OA
1MA
1LA
1KA
1JA
0HA
0GA
0@A
1>A
1=A
1$B
1"B
0{A
0yA
1wA
1vA
0uA
0VD
0TD
1ED
1DD
1CD
0>D
0:D
06D
1QE
1PE
1OE
0NE
0LE
0JE
1HE
0DE
1CE
0BE
1@E
0?E
1>E
1;E
09E
07E
05E
04E
13E
12E
01E
0/E
1-E
1,E
0+E
0*E
0)E
1zE
1vE
0uE
1rE
0oE
0lE
0jE
1hE
0gE
1eE
1dE
1aE
1`E
0_E
1]E
1[E
1VE
0cP
0[P
0YP
0OP
1NP
0KP
1IP
0HP
1>P
0<P
07P
06P
04P
02P
1BO
0AO
0@O
1:O
19O
18O
15O
02O
01O
00O
0/O
1.O
1-O
0,O
0+O
0*O
0)O
1&O
0$O
1"O
1!O
1{N
0zN
0yN
1wN
0vN
0uN
1qN
1pN
0oN
0nN
1jN
1iN
0hN
0gN
0fN
0eN
1dN
1cN
1bN
1#P
1qO
1oO
1jO
1iO
0fO
1dO
0bO
0aO
0]O
1[O
1WO
1VO
1UO
1TO
1QO
1PO
0OO
1HO
1AO
09O
17O
0-O
1,O
1)O
0'O
0&O
1zN
1xN
1sN
1rN
0pN
1nN
0#P
0wO
0iO
1gO
0ZO
0UO
0TO
0PO
0PE
1NE
1?E
0>E
1=E
08E
14E
10E
0zE
1jE
0`E
0\E
1bA
0_A
0^A
0\A
0XA
0WA
0VA
1SA
1GA
10B
1(B
0$B
0vA
1k=
0b=
1S=
08>
0~=
#75600
b10001001001100101101011000010010 d
b1000111111011001101101110001111 e
0"
1&Y
0%Y
0$Y
0#Y
1"Y
1!Y
1|X
0zX
1xX
0vX
1uX
1tX
0sX
1rX
1mX
0lX
0kX
0jX
1iX
0hX
1r!
0q!
0p!
0o!
1n!
1m!
1j!
0h!
1f!
0d!
1c!
1b!
0a!
1`!
1[!
0Z!
0Y!
0X!
1W!
0V!
0gX
1fX
0eX
1cX
0bX
0aX
0`X
0_X
0ZX
0WX
0UX
0TX
1SX
0PX
1OX
0NX
1LX
0KX
0JX
0IX
1HX
0G!
1E!
1D!
0C!
0B!
0A!
0?!
1>!
0=!
1<!
19!
18!
15!
13!
1.!
0,!
1+!
1*!
1$!
0~
0}
1|
1{
0y
1x
0w
0v
1u
1t
1r
0p
0o
1n
0m
1l
1k
1j
1i
0h
0T!
1o(
0n(
0m(
0l(
1k(
1j(
1g(
0e(
1c(
0a(
1`(
1_(
0^(
1](
1X(
0W(
0V(
0U(
1T(
0S(
07"
16"
05"
13"
02"
01"
00"
0/"
0*"
0'"
0%"
0$"
1#"
0~!
1}!
0|!
1z!
0y!
0x!
0w!
1v!
b1 yQ
b0 vQ
b1 sQ
b0 mQ
b0 pQ
b1 dQ
b0 ^Q
b1 aQ
b1 XQ
b0 RQ
b1 LQ
1PQ
0YQ
1\Q
0bQ
0eQ
0kQ
b101110000001001100100100011100001 KQ
b1000111111011001101101110001111 NQ
b1000111111011001101101110001111 QQ
b101110000001001100100100011100001 WQ
b10001111110110011011011100011110 ZQ
b1000111111011001101101110001111 ]Q
b110111000000100110010010001110000 `Q
b110111000000100110010010001110000 cQ
b1000111111011001101101110001111 fQ
b110111000000100110010010001110000 iQ
b1000111111011001101101110001111 lQ
b1000111111011001101101110001111 oQ
b101110000001001100100100011100001 rQ
b1000111111011001101101110001111 uQ
b101110000001001100100100011100001 xQ
1$)
0!)
1~(
0|(
0{(
0y(
1q'
0p'
0o'
0n'
0g'
1f'
0d'
0b'
1`'
0Z'
0Y'
0X'
0W'
1P'
1O'
1N'
1G'
0F'
1D'
1B'
0@'
1:'
19'
18'
17'
0.'
0-'
0+'
1('
0&'
1$'
0#'
0"'
1{&
0y&
1x&
0w&
0v&
0u&
0t&
0r&
1o&
0n&
1l&
1k&
1j&
1c&
0b&
1`&
1^&
0\&
1V&
1U&
1T&
1S&
1K&
1J&
1I&
1B&
0A&
1?&
1=&
0;&
15&
14&
13&
12&
0'&
1&&
1%&
1$&
0#&
0"&
0}%
1{%
0y%
1w%
0v%
0u%
1t%
0s%
0n%
1m%
1l%
1k%
0j%
1i%
1h%
1g%
1f%
1e%
1d%
1`%
1_%
1^%
1\%
1[%
1Y%
1X%
1U%
1T%
1R%
1Q%
1P%
1O%
1N%
1M%
1I%
1B%
1A%
1@%
1<%
19%
16%
15%
12%
1+%
1*%
1)%
1'%
1&%
1!%
1~$
1}$
1y$
1v$
1s$
1r$
1o$
1h$
1g$
1f$
1d$
1c$
1b$
1a$
1`$
1Y$
0X$
1V$
1T$
0R$
1L$
1K$
1J$
1I$
1=$
0<$
0;$
0:$
19$
18$
15$
03$
11$
0/$
1.$
1-$
0,$
1+$
1&$
0%$
0$$
0#$
1"$
0!$
1~#
1y#
1x#
1w#
1s#
1p#
1m#
1l#
1i#
1b#
1a#
1`#
1^#
1;#
1:#
19#
08#
15#
1.#
1-#
0,#
0+#
1*#
0(#
1'#
1%#
1$#
1##
1"#
0!#
1|"
0{"
1v"
0u"
0t"
0s"
1r"
1q"
1n"
0l"
1j"
0h"
1g"
1f"
0e"
1d"
1_"
0^"
0]"
0\"
1["
0Z"
0Y"
0W"
0V"
0T"
1Q"
0O"
1M"
0L"
0K"
1F"
0D"
1C"
0B"
0A"
0@"
0?"
0="
1:"
09"
14(
08(
1<(
1B(
0@(
1D(
0L(
0J(
1N(
0P(
1R(
1m8
0U,
0l)
0k)
0i)
1f)
0d)
1b)
0a)
0`)
1[)
0Y)
1X)
0W)
0V)
0U)
0T)
0R)
1O)
0N)
1,,
1+,
1*,
0),
1&,
1}+
1|+
0{+
0z+
1y+
0w+
1v+
1t+
1s+
1r+
1q+
0p+
1m+
0l+
1Q/
1P/
1O/
1H/
0G/
1E/
1C/
0A/
1;/
1:/
19/
18/
1Q2
1O2
1N2
1M2
1L2
1H2
1G2
1F2
1D2
1C2
1A2
1@2
1=2
1<2
1:2
192
182
172
162
152
112
1'5
1&5
1%5
1|4
0{4
1y4
1w4
0u4
1o4
1n4
1m4
1l4
0O5
1M5
1L5
1K5
1D5
0C5
1A5
1?5
0=5
175
165
155
145
0u5
0r5
0q5
0o5
1l5
0j5
1h5
0g5
0f5
1a5
0_5
1^5
0]5
0\5
0[5
0Z5
0X5
1U5
0T5
1%8
1#8
1"8
1!8
1x7
0w7
1u7
1s7
0q7
1k7
1j7
1i7
1h7
0I8
1G8
0F8
0E8
0D8
0=8
1<8
0:8
088
168
008
0/8
0.8
0-8
0r2
1q2
1p2
1o2
0n2
0m2
0j2
1h2
0f2
1d2
0c2
0b2
1a2
0`2
0[2
1Z2
1Y2
1X2
0W2
1V2
1U2
0T2
1+2
1%2
1$2
1#2
1}1
1z1
1w1
1v1
1s1
1l1
1k1
1j1
1h1
1g1
0f1
0y/
1s/
1r/
1q/
1m/
1j/
1g/
1f/
1c/
1\/
1[/
1Z/
1X/
1W/
0V/
1-/
1'/
0&/
0%/
0$/
1#/
1"/
1}.
0{.
1y.
0w.
1v.
1u.
0t.
1s.
1n.
0m.
0l.
0k.
1j.
0i.
1h.
1y,
1t,
1s,
1r,
1n,
1k,
1h,
1g,
1d,
1],
1\,
1[,
1Y,
0X,
13*
1.*
0-*
0,*
0+*
1**
1)*
1&*
0$*
1"*
0~)
1})
1|)
0{)
1z)
1u)
0t)
0s)
0r)
1q)
0p)
0o)
1n)
127
017
007
0/7
1.7
0-7
1+7
1*7
0)7
1&7
0$7
1#7
1"7
0!7
0z6
0y6
1x6
1u6
0t6
0r6
1o6
1n6
1Y7
1X7
1W7
0V7
0S7
1P7
0N7
1M7
1L7
0K7
0J7
1E7
1D7
1C7
1B7
0?7
087
174
154
134
124
1/4
0.4
1-4
1+4
0)4
0'4
0&4
1$4
0"4
0}3
1y3
1v3
0u3
1s3
0q3
0p3
1o3
0n3
1Y4
1X4
1T4
1S4
1P4
1O4
1M4
1L4
1I4
1H4
1E4
1B4
1A4
1>4
1=4
1:4
191
041
121
011
001
1-1
1,1
0)1
0&1
1$1
1!1
0|0
0{0
1y0
0x0
0w0
0r0
1q0
0p0
1\1
1[1
0Z1
1W1
1V1
1Q1
1O1
1N1
0M1
1K1
1G1
1F1
1E1
1D1
0C1
1@1
1>1
1<1
0A+
0@+
1?+
1=+
0<+
1;+
09+
17+
06+
05+
02+
00+
1/+
0.+
1)+
1(+
1&+
0%+
1$+
0!+
1~*
1}*
1|*
1e+
0c+
0a+
1`+
0_+
1Z+
1T+
1P+
0O+
0M+
0L+
0J+
1I+
0H+
0F+
1E+
0D+
0C+
19.
18.
17.
16.
12.
00.
1/.
0..
1+.
0).
0(.
0%.
0#.
1".
1!.
1}-
0|-
1y-
0x-
1w-
0v-
1u-
1s-
0r-
0a.
1X.
1V.
1R.
1O.
1L.
1K.
1H.
1@.
1':
1$:
1#:
1":
0!:
0~9
0z9
1y9
1v9
0u9
1t9
0s9
0r9
0p9
0m9
0l9
0k9
0i9
0h9
1g9
1I:
0H:
1B:
0A:
1=:
0<:
18:
15:
14:
13:
0/:
#77400
1"
1T!
b111001101111100101010010011011011100 N:
b100010000001000100100100000100001 O:
b111010100010110001000010101011001111100 P:
b100000001001100100100010100000000000 Q:
b100000001000101011000100111100010001001 R:
b10111000111110110011011001110001110000 S:
b100110010011010010010000011010100110101 T:
b10011001100100110011011001100011000000 U:
b111000101101000111011001110111010001101 V:
b110000011111100100110011100001110000 W:
b101101001000100000101011010000111101 X:
b1010100010111011101010100111000010000 Y:
b101011011000101110100010011110100101110011 "F
b10000001001000100000001000000000 #F
b1011101110101011111001001000001110100001001000 $F
b100000000100100100000001000000000 %F
b10001110101110000001010111010000100101110101 &F
b101001010001101110101000100111001000000000 'F
b100011111010011100110101011001011010010011010011010010 xK
b100010001010100111000101101100100000000000 yK
b1110001000100001101111001100101010011111010100000000000 zK
b1000101001100010000010010100000100000000000000000000 {K
b1110000111101001110001101111111101001100101000001111101010010110 HQ
b100000000100001100010000000010010010000101000000000000000000 IQ
b1101111010011111001011100101100001110111000111101111101000001110 P!
b1110000101110100110110011101000001001101000010100011010101110011 Q!
b10011011110001011010010110110000110111001101100010011010010 R!
b1111000111110010001010010000000001110000110010001111101010010110 S!
b10001001001100101101011000010010 H!
b1110010101011111111011111100101 J!
b11100010111101111000010011000101 L!
b1111100111111011110100111111001 N!
b1000111111011001101101110001111 I!
b10111011110100100111001001110111 K!
b11010101000100111101001010101010 M!
b11100011001101110010010011000110 O!
1iY
1dY
0bY
1aY
1]Y
1\Y
0[Y
0ZY
0WY
1VY
0TY
0SY
0RY
1QY
0PY
1NY
1KY
0JY
0IY
0GY
0FY
1EY
0DY
1CY
1BY
0?Y
1=Y
0<Y
1;Y
1:Y
08Y
06Y
14Y
02Y
11Y
0/Y
1,Y
1+Y
1*Y
1b
0`
1Z
1X
1W
1V
0R
0Q
0O
1M
0K
0J
0I
0H
1F
1E
0B
0A
0=
1;
0:
09
18
05
03
1.
1-
1+
1'
1%
1$
0GN
0FN
1=N
05N
12N
0/N
1.N
1-N
0,N
1*N
1(N
0&N
1$N
0lM
1kM
1iM
1gM
1fM
1eM
1cM
0_M
1^M
0]M
1YM
1UM
1PM
0MM
0HM
0GM
1FM
0DM
13M
01M
1/M
0.M
1-M
1,M
1*M
0)M
0'M
1&M
1%M
1}L
0|L
0xL
0[L
1WL
0TL
1SL
0RL
1ML
0LL
0KL
0IL
0DL
1BL
1=L
01L
10L
1-L
1,L
0*L
1RJ
0QJ
1NJ
1JJ
0HJ
1AJ
1@J
1=J
0;J
0:J
19J
08J
17J
12J
1#J
1!J
0|I
0zI
1xI
0tI
1sI
0rI
1pI
1mI
1kI
0iI
0hI
0gI
0eI
1cI
1bI
0aI
1`I
0_I
1]I
1\I
0[I
0ZI
0YI
1NI
0JI
0HI
1FI
1@I
0=I
0;I
09I
17I
05I
03I
0-I
0aG
1`G
0_G
0^G
0\G
1[G
0ZG
1YG
1WG
0VG
0UG
0TG
0SG
0OG
0MG
1KG
1JG
1IG
1HG
0FG
0>G
1<G
1;G
0)G
0&G
1%G
1!G
0}F
1|F
1uF
0tF
0pF
0lF
1^F
1YF
0WF
1VF
0RF
1QF
1NF
0MF
0LF
0JF
0IF
1GF
0FF
1CF
0BF
0@F
0?F
1=F
0;F
1:F
08F
17F
15F
1"D
0!D
1yC
0xC
1tC
0sC
1oC
1lC
1kC
1jC
0fC
1YC
1VC
1UC
1TC
0SC
0RC
0NC
1MC
1JC
0IC
1HC
0GC
0FC
0DC
0AC
0@C
0?C
0=C
0<C
1;C
1.C
1-C
1,C
0+C
0(C
1%C
0#C
1"C
1!C
0~B
0}B
1xB
1wB
1vB
1uB
0rB
0kB
1bB
0aB
0`B
0_B
1^B
0]B
1[B
1ZB
0YB
1VB
0TB
1SB
1RB
0QB
0LB
0KB
1JB
1GB
0FB
0DB
1AB
1@B
1,@
1+@
1'@
1&@
1#@
1"@
1~?
1}?
1z?
1y?
1v?
1s?
1r?
1o?
1n?
1k?
1b?
1`?
1^?
1]?
1Z?
0Y?
1X?
1V?
0T?
0R?
0Q?
1O?
0M?
0J?
1F?
1C?
0B?
1@?
0>?
0=?
1<?
0;?
13?
12?
01?
1.?
1-?
1(?
1&?
1%?
0$?
1"?
1|>
1{>
1z>
1y>
0x>
1u>
1s>
1q>
1h>
0c>
1a>
0`>
0_>
1\>
1[>
0X>
0U>
1S>
1P>
0M>
0L>
1J>
0I>
0H>
0C>
1B>
0A>
0D<
1;<
19<
15<
12<
1/<
1.<
1+<
1#<
1x;
1w;
1v;
1u;
1q;
0o;
1n;
0m;
1j;
0h;
0g;
0d;
0b;
1a;
1`;
1^;
0];
1Z;
0Y;
1X;
0W;
1V;
1T;
0S;
1P;
0N;
0L;
1K;
0J;
1E;
1?;
1;;
0:;
08;
07;
05;
14;
03;
01;
10;
0/;
0.;
0&;
0%;
1$;
1";
0!;
1~:
0|:
1z:
0y:
0x:
0u:
0s:
1r:
0q:
1l:
1k:
1i:
0h:
1g:
0d:
1c:
1b:
1a:
0NR
1LR
1KR
1JR
1GR
0FR
1DR
0CR
1?R
0=R
0;R
18R
17R
16R
14R
13R
10R
1?=
1==
0<=
1;=
17=
16=
04=
02=
1/=
0-=
1)=
1&=
0%=
1$=
0!=
1~<
1}<
0|<
1uR
1sR
1rR
1nR
0lR
0jR
0iR
1gR
0dR
0bR
0aR
1]R
0ZR
1WR
0VR
1UR
0TR
1QR
0PR
1+>
1)>
1%>
1|=
1y=
1q=
1vS
1qS
1pS
0mS
0kS
0iS
1fS
0eS
1bS
1_S
0^S
1YS
0VS
1TS
1RS
0QS
0OS
19A
04A
12A
01A
1.A
1-A
1+A
0)A
0#A
0|@
1y@
0x@
1r@
1q@
1AT
1?T
1=T
1<T
1:T
08T
17T
04T
03T
1-T
0,T
1*T
0&T
1%T
1#T
0!T
0|S
0{S
0zS
0xS
1'B
1&B
1#B
1~A
1}A
1zA
1sA
1oA
1kA
1BU
0AU
1;U
19U
07U
16U
05U
1)U
1'U
0$U
0!U
1~T
1}T
1$E
1!E
1~D
0}D
1|D
1{D
1zD
0yD
1vD
0tD
1sD
0qD
0oD
1nD
0mD
0lD
1jD
1gD
0fD
0eD
0bD
1aD
1`D
1kU
1hU
1gU
0dU
1`U
1^U
0\U
0[U
1XU
1VU
1UU
0SU
0PU
0OU
1NU
1MU
0LU
0sE
1mE
1cE
1_E
1^E
1GH
1BH
0@H
1?H
0;H
18H
15H
04H
01H
0/H
1-H
0+H
0)H
0'H
1&H
0~G
0}G
0uG
1sG
1rG
0oH
0mH
0lH
1kH
0jH
1hH
1gH
0fH
0dH
0_H
1^H
0]H
1ZH
1WH
17K
0/K
0.K
1,K
1+K
1)K
1'K
1%K
0#K
1!K
1~J
0}J
0|J
0{J
0zJ
1yJ
1uJ
1sJ
0nJ
1mJ
1lJ
1kJ
0jJ
1fK
0cK
0]K
0[K
1ZK
0XK
1VK
1TK
0RK
0NK
0JK
1IK
0HK
1GK
0DK
0"W
1|V
0yV
1xV
0wV
0vV
0tV
0oV
0nV
0mV
1lV
1jV
1hV
0gV
0aV
0]V
0VV
1UV
1RV
1QV
0OV
1AQ
1=Q
17Q
06Q
04Q
13Q
1.Q
1+Q
1'Q
1&Q
1{P
1xP
1vP
1uP
1tP
0QW
1PW
1NW
1LW
1KW
1IW
1HW
0DW
1CW
0BW
1@W
0>W
1:W
18W
11W
10W
1/W
0,W
0'W
1_O
0QO
1OO
1JO
0HO
1^P
1ZP
1TP
0SP
0QP
1PP
1KP
1HP
1DP
1CP
1:P
17P
15P
14P
13P
0DX
1@X
0=X
1<X
0;X
0:X
08X
01X
0-X
0,X
0*X
0&X
0$X
1"X
0!X
0~W
0zW
0wW
0tW
1sW
1pW
0oW
0lW
0gW
0AQ
0=Q
1;Q
14Q
03Q
12Q
1-Q
0&Q
0yP
0tP
1UD
1RD
1QD
0PD
1OD
1ND
1MD
0LD
1ID
0GD
1FD
0DD
0BD
1AD
0@D
0?D
1=D
1:D
09D
08D
05D
14D
13D
1<V
0;V
09V
06V
13V
02V
01V
10V
0/V
0.V
0,V
0*V
1)V
0&V
1$V
0{U
0zU
0wU
0$E
1wD
0vD
0uD
0gD
0dD
0`D
1g@
0b@
1`@
0_@
1\@
1[@
1Y@
0W@
0Q@
0L@
1I@
0H@
1B@
1A@
1vT
1qT
1nT
0mT
1lT
0gT
0eT
1cT
0_T
0^T
1\T
1[T
0VT
0UT
0QT
0PT
0OT
0MT
0LT
0KT
0IT
09A
13A
1,A
1)A
1(A
1!A
1u@
0r@
1q<
1o<
0n<
1m<
1i<
1h<
0f<
0d<
1a<
0_<
1[<
1X<
0W<
1V<
0S<
1R<
1Q<
0P<
0FS
1DS
1CS
1@S
1>S
1<S
19S
16S
05S
14S
03S
01S
10S
0,S
1+S
1*S
1(S
0'S
0$S
1#S
1"S
0!S
1|R
0{R
0?=
0>=
09=
07=
06=
0)=
0'=
0q<
0p<
0k<
0i<
0h<
0[<
0Y<
0l=
1j=
0g=
1e=
0d=
1b=
0a=
1`=
0_=
0^=
1[=
1Z=
1V=
0S=
0R=
0Q=
0O=
1M=
0K=
0G=
1D=
0C=
16>
14>
11>
1.>
1,>
0)>
0(>
0$>
1~=
1}=
1{=
0x=
1t=
0g@
1a@
1Z@
1W@
1V@
1O@
1E@
0B@
1hA
1gA
1cA
0bA
1^A
1\A
0[A
1UA
0PA
1NA
0MA
0LA
0IA
0GA
0CA
0?A
0>A
0=A
0;A
11B
00B
1,B
0(B
0&B
0}A
1|A
1xA
0wA
1vA
1rA
1nA
0UD
1JD
0ID
0HD
0:D
07D
03D
1PE
0ME
1LE
0KE
1IE
0HE
1EE
1DE
1BE
0AE
0=E
1<E
0;E
19E
18E
17E
04E
03E
02E
11E
00E
1/E
0.E
1wE
0vE
1tE
1sE
0rE
0qE
1oE
1iE
0hE
1gE
0eE
0dE
1`E
0]E
1\E
0[E
1ZE
0^P
0ZP
1XP
1QP
0PP
1OP
1JP
0CP
08P
03P
0AO
1=O
0<O
0:O
19O
07O
05O
12O
11O
1/O
1*O
1'O
1&O
0#O
0"O
0}N
0|N
0{N
0wN
1vN
1tN
0sN
1oN
1mN
0lN
0iN
0dN
1|O
0qO
0oO
0jO
0gO
1bO
1]O
0VO
1UO
1RO
0OO
1FO
1<O
08O
06O
0/O
0.O
1-O
0(O
0!O
0tN
0oN
0|O
1vO
1oO
1hO
0OE
0DE
0CE
0BE
14E
01E
0-E
1pE
0`E
0gA
1aA
0ZA
1WA
1VA
1OA
0EA
0BA
1+B
1tA
1i=
0h=
1c=
1a=
0`=
1S=
1Q=
06>
00>
0.>
0~=
0|=
#79200
b1111001001100000110100111110010 d
b11100111011101101001011011001110 e
0"
0)Y
1#Y
0!Y
1}X
0|X
0yX
1vX
0tX
1sX
0pX
1jX
1hX
0u!
1o!
0m!
1k!
0j!
0g!
1d!
0b!
1a!
0^!
1X!
1V!
1bX
1aX
1`X
1_X
0^X
0]X
1\X
0[X
1ZX
0XX
0VX
1KX
1JX
1IX
0HX
0F!
1C!
1B!
1@!
0>!
1=!
0;!
0:!
09!
08!
17!
06!
04!
10!
0/!
0*!
0)!
1%!
1}
0|
0{
1w
0u
0s
0r
0q
1p
1o
0n
0l
0j
1h
0T!
0r(
1l(
0j(
1h(
0g(
0d(
1a(
0_(
1^(
0[(
1U(
1S(
12"
11"
10"
1/"
0."
0-"
1,"
0+"
1*"
0("
0&"
1y!
1x!
1w!
0v!
b0 yQ
b0 dQ
b0 aQ
b1 ^Q
b1 [Q
b0 XQ
b1 RQ
1MQ
0PQ
1eQ
1kQ
0nQ
0qQ
1tQ
b110001000100101101001001100011 KQ
b111100111011101101001011011001110 NQ
b11000100010010110100100110001 QQ
b111001110111011010010110110011100 WQ
b110001000100101101001001100011 ZQ
b11000100010010110100100110001 ]Q
b111001110111011010010110110011100 `Q
b0 cQ
b0 fQ
b11000100010010110100100110001 iQ
b111100111011101101001011011001110 lQ
b111100111011101101001011011001110 oQ
b110001000100101101001001100011 rQ
b0 uQ
b111001110111011010010110110011100 xQ
1%)
0$)
1{(
1y(
0x(
0w(
1v(
0q'
1o'
1n'
1m'
0l'
0k'
1i'
1g'
1d'
0c'
1a'
0`'
1^'
1['
1Z'
1X'
1W'
1V'
0U'
0T'
1R'
0P'
0O'
0N'
0M'
0I'
0H'
0G'
0E'
0D'
0B'
0A'
0>'
0='
0;'
0:'
09'
08'
07'
06'
02'
1.'
0('
1&'
0$'
1#'
1~&
0{&
1y&
0x&
1u&
0o&
0m&
0l&
1f&
0d&
1b&
0a&
0^&
1[&
0Y&
1X&
0U&
1O&
1M&
1L&
0K&
1E&
0C&
1A&
0@&
0=&
1:&
08&
17&
04&
1.&
1,&
1+&
1*&
0$&
1"&
0~%
1}%
1z%
0w%
1u%
0t%
1q%
0k%
0i%
0h%
0g%
0f%
0e%
0d%
0`%
0_%
0^%
0\%
0[%
0Y%
0X%
0U%
0T%
0R%
0Q%
0P%
0O%
0N%
0M%
0I%
0B%
0A%
0@%
0<%
09%
06%
05%
02%
0+%
0*%
0)%
0'%
0&%
1#%
1"%
0~$
0}$
1|$
1{$
1x$
0r$
1q$
1p$
0o$
1n$
1m$
1l$
1j$
1i$
0g$
0f$
1e$
0a$
0`$
0_$
1^$
1]$
0[$
0Y$
0V$
1U$
0S$
1R$
0P$
0M$
0L$
0J$
0I$
0H$
1G$
1F$
0D$
1A$
0?$
0>$
0=$
1<$
1;$
09$
07$
04$
13$
01$
10$
0.$
0+$
0*$
0($
0'$
0&$
1%$
1$$
0"$
0~#
1|#
1{#
1z#
0y#
0x#
1v#
1t#
1q#
0p#
1n#
0m#
1k#
1h#
1g#
1e#
1d#
1c#
0b#
0a#
1_#
0;#
0:#
09#
18#
17#
05#
03#
00#
1/#
0-#
1,#
0*#
0'#
0&#
0$#
0##
0"#
1!#
1~"
0|"
0y"
1s"
0q"
1o"
0n"
0k"
1h"
0f"
1e"
0b"
1\"
1Z"
1Y"
1W"
0Q"
1O"
0M"
1L"
1I"
0F"
1D"
0C"
1@"
0:"
08"
18(
0<(
1>(
1@(
0B(
0D(
0R(
0m8
1U,
0,,
0+,
0*,
1),
1(,
0&,
0$,
0!,
1~+
0|+
1{+
0y+
0v+
0u+
0s+
0r+
0q+
1p+
1o+
0m+
0y,
1w,
1v,
1u,
0t,
0s,
1q,
1o,
1l,
0k,
1i,
0h,
1f,
1c,
1b,
1`,
1_,
1^,
0],
0\,
1Z,
0-/
1+/
0)/
0(/
0'/
1&/
1%/
0#/
0!/
0|.
1{.
0y.
1x.
0v.
0s.
0r.
0p.
0o.
0n.
1m.
1l.
0j.
1S/
0P/
0O/
0N/
1M/
1L/
0J/
0H/
0E/
1D/
0B/
1A/
0?/
0</
0;/
09/
08/
07/
16/
15/
03/
1y/
1u/
1t/
0r/
0q/
1p/
1o/
1l/
0f/
1e/
1d/
0c/
1b/
1a/
1`/
1^/
1]/
0[/
0Z/
1Y/
0Q2
0O2
0N2
0M2
0L2
0H2
0G2
0F2
0D2
0C2
0A2
0@2
0=2
0<2
0:2
092
082
072
062
052
012
0#8
0"8
0!8
0~7
0z7
0y7
0x7
0v7
0u7
0s7
0r7
0o7
0n7
0l7
0k7
0j7
0i7
0h7
0g7
0c7
0G8
1E8
1D8
1C8
0B8
0A8
1?8
1=8
1:8
098
178
068
148
118
108
1.8
1-8
1,8
0+8
0*8
1(8
1r5
0l5
1j5
0h5
1g5
1d5
0a5
1_5
0^5
1[5
0U5
0S5
1R5
0M5
1G5
0E5
1C5
0B5
0?5
1<5
0:5
195
065
105
1.5
1-5
0,5
0'5
1!5
0}4
1{4
0z4
0w4
1t4
0r4
1q4
0n4
1h4
1f4
1e4
0d4
1u2
0o2
1m2
0k2
1j2
1g2
0d2
1b2
0a2
1^2
0X2
0V2
0U2
1T2
0+2
0%2
0$2
0#2
0}1
0z1
0w1
0v1
0s1
0l1
0k1
0j1
0h1
0g1
1f1
01*
1+*
0)*
1'*
0&*
0#*
1~)
0|)
1{)
0x)
1r)
1p)
1o)
0n)
1l)
0f)
1d)
0b)
1a)
1^)
0[)
1Y)
0X)
1U)
0O)
0M)
0L)
0K)
1J)
1@+
0?+
0:+
19+
08+
07+
16+
04+
12+
01+
0/+
1.+
0-+
1++
0)+
0(+
0#+
1"+
1!+
1\+
0Z+
1Y+
1Q+
0P+
1M+
0E+
037
117
0.7
1-7
0'7
1%7
1$7
0"7
0~6
0}6
0|6
1z6
1y6
0u6
1t6
1q6
0n6
0m6
1l6
0Y7
1V7
0P7
1O7
0M7
0L7
1J7
1H7
1G7
0D7
0B7
1?7
1<7
074
054
034
024
114
0/4
1,4
0+4
0*4
1)4
1&4
1#4
0z3
0y3
1x3
0v3
1t3
1p3
0o3
1n3
0Y4
0X4
0T4
0S4
0P4
0O4
0M4
0L4
0I4
0H4
0E4
0B4
0A4
0>4
0=4
0:4
091
111
1/1
0+1
1*1
1'1
1%1
0$1
0#1
1"1
1~0
1{0
1z0
1x0
1v0
1t0
1s0
1_1
0\1
0[1
1Y1
1X1
0W1
0V1
0U1
1S1
0R1
1P1
0O1
0J1
0H1
0G1
0E1
0D1
1B1
1A1
0@1
0?1
0>1
09.
08.
07.
06.
14.
13.
01.
0/.
1,.
0+.
1*.
1).
1(.
1%.
1#.
0".
0!.
1~-
1{-
1z-
1x-
0w-
1v-
0t-
1a.
1Y.
0X.
1S.
0R.
0O.
0L.
0K.
1J.
0H.
1F.
0@.
1>.
0%:
0$:
0#:
0":
1!:
1~9
1}9
1z9
0y9
0x9
1u9
1s9
1m9
1l9
1i9
1h9
0g9
1f9
0d9
0b9
0I:
0D:
0C:
0B:
1A:
0=:
0;:
08:
05:
04:
01:
1/:
0-:
1*:
#81000
1"
1T!
b111110101100110010001000100101011010 N:
b10001000100100101001000100001 O:
b101101111011001011011101100001111000000 P:
b10000000100010000000010010010000000100 Q:
b101101011110111100101101011110110001000 R:
b10000110001000010010110100001100010100 S:
b1010111000100010010110100100110001000000 T:
b0 U:
b1001010110101110000001111010111100011001 V:
b111001010101111110000101100011100000 W:
b110111011100001111000110111000001 X:
b1110001000100010100000101000000000000 Y:
b11001010010001010110011111000111011001110 "F
b100100001010101000100000110000100100000 #F
b1000000001100110001011101001110010101001 $F
b100110011101010101010110101000110000100000000 %F
b10001001000010011100100110000100010010101101 &F
b101010101101110011011001111001100100000000 'F
b101110111010000100111000001100001001011010010101110011 xK
b101011000100100010110010000100100000000000 yK
b1101110000110101110000111001111111110011010101000000000 zK
b1010001000000101000100000000000100000000000000000 {K
b1100000011011001100010101000100001110110110001101000010011010010 HQ
b10001000000010010100010101001010001000000100000010000000000000 IQ
b1111010001100010011010010101110000010110100101010000110010111100 P!
b1101111010011111001011100101100001110111000111101111101000001110 Q!
b1110000101110100110110011101000001001101000010100011010101110011 R!
b10011011110001011010010110110000110111001101100010011010010 S!
b1111001001100000110100111110010 H!
b10001001001100101101011000010010 J!
b1110010101011111111011111100101 L!
b11100010111101111000010011000101 N!
b11100111011101101001011011001110 I!
b1000111111011001101101110001111 K!
b10111011110100100111001001110111 M!
b11010101000100111101001010101010 O!
0iY
1gY
1fY
0eY
0dY
0cY
0aY
1`Y
0_Y
1^Y
1[Y
1ZY
1WY
1UY
1PY
0NY
1MY
1LY
1FY
0BY
0AY
1@Y
1?Y
0=Y
1<Y
0;Y
0:Y
19Y
18Y
16Y
04Y
03Y
12Y
01Y
10Y
1/Y
1.Y
1-Y
0,Y
0a
1]
0Z
1Y
0X
0W
0V
1R
1Q
0P
1N
1J
1I
0G
0F
0E
1D
1C
1A
1@
1>
19
11
10
0.
0+
1)
0'
0&
0%
0$
1FN
0CN
0=N
0;N
1:N
08N
16N
14N
02N
0.N
0*N
1)N
0(N
1'N
0$N
1mM
0eM
0dM
1bM
1aM
1_M
1]M
1[M
0YM
1WM
1VM
0UM
0TM
0SM
0RM
1QM
1MM
1KM
0FM
1EM
1DM
1CM
0BM
0/M
0-M
0,M
1+M
0*M
1(M
1'M
0&M
0$M
0}L
1|L
0{L
1xL
1uL
1]L
1XL
0VL
1UL
0QL
1NL
1KL
0JL
0GL
0EL
1CL
0AL
0?L
0=L
1<L
06L
05L
0-L
1+L
1*L
1SJ
0RJ
1PJ
0NJ
0MJ
1LJ
1KJ
1IJ
1EJ
0DJ
1CJ
0AJ
0@J
1?J
1;J
1:J
09J
18J
07J
16J
1"J
0!J
0}I
1|I
0{I
1yI
0xI
1uI
0sI
0qI
0mI
1lI
0kI
1iI
1hI
1gI
0cI
0bI
0`I
1_I
0^I
0]I
1OI
0NI
1JI
1II
0FI
1EI
1AI
1>I
1<I
1:I
18I
07I
16I
14I
13I
12I
1/I
1.I
1+I
1fG
1aG
0`G
1_G
1\G
1ZG
0YG
0XG
1UG
1TG
1SG
0NG
1MG
1LG
0KG
0JG
0GG
0EG
0CG
0AG
0@G
0=G
0<G
0;G
09G
11G
1.G
0-G
1)G
1(G
0%G
1"G
0!G
1zF
1xF
1vF
0uF
1qF
1nF
0^F
1\F
1[F
0ZF
0YF
1WF
0VF
1UF
1TF
0QF
0PF
1MF
1LF
1HF
0DF
0AF
1?F
0=F
09F
16F
05F
0"D
0{C
0zC
0yC
1xC
0tC
0rC
0oC
0lC
0kC
0hC
1fC
0dC
1aC
0WC
0VC
0UC
0TC
1SC
1RC
1QC
1NC
0MC
0LC
1IC
1GC
1AC
1@C
1=C
1<C
0;C
1:C
08C
06C
0.C
1+C
0%C
1$C
0"C
0!C
1}B
1{B
1zB
0wB
0uB
1rB
1oB
0cB
1aB
0^B
1]B
0WB
1UB
1TB
0RB
0PB
0OB
0NB
1LB
1KB
0GB
1FB
1CB
0@B
0?B
1>B
0,@
0+@
0'@
0&@
0#@
0"@
0~?
0}?
0z?
0y?
0v?
0s?
0r?
0o?
0n?
0k?
0b?
0`?
0^?
0]?
1\?
0Z?
1W?
0V?
0U?
1T?
1Q?
1N?
0G?
0F?
1E?
0C?
1A?
1=?
0<?
1;?
16?
03?
02?
10?
1/?
0.?
0-?
0,?
1*?
0)?
1'?
0&?
0!?
0}>
0|>
0z>
0y>
1w>
1v>
0u>
0t>
0s>
0h>
1`>
1^>
0Z>
1Y>
1V>
1T>
0S>
0R>
1Q>
1O>
1L>
1K>
1I>
1G>
1E>
1D>
1D<
1<<
0;<
16<
05<
02<
0/<
0.<
1-<
0+<
1)<
0#<
1!<
0x;
0w;
0v;
0u;
1s;
1r;
0p;
0n;
1k;
0j;
1i;
1h;
1g;
1d;
1b;
0a;
0`;
1_;
1\;
1[;
1Y;
0X;
1W;
0U;
1G;
0E;
1D;
1<;
0;;
18;
00;
1%;
0$;
0}:
1|:
0{:
0z:
1y:
0w:
1u:
0t:
0r:
1q:
0p:
1n:
0l:
0k:
0f:
1e:
1d:
0MR
0LR
0GR
1FR
0ER
1CR
0BR
0?R
0>R
1<R
1;R
0:R
19R
06R
00R
1/R
1.R
1-R
0==
0:=
19=
18=
17=
16=
05=
0/=
1.=
1-=
1)=
1'=
0&=
1"=
1!=
1|<
0uR
0sR
0rR
1pR
1oR
0mR
1lR
1hR
0gR
1dR
1bR
1aR
1\R
1[R
1XR
1VR
0UR
1TR
1SR
0RR
0QR
0+>
1&>
0%>
0}=
1w=
0q=
0vS
0sS
0pS
1oS
1nS
1mS
1kS
1jS
1iS
0hS
0fS
0cS
0bS
0aS
0`S
0_S
1^S
1]S
1\S
0[S
0ZS
1XS
1WS
1VS
0TS
03A
11A
1/A
0+A
1*A
1'A
0&A
1%A
1"A
1~@
1x@
1v@
0u@
1t@
0AT
0?T
0=T
0<T
1;T
0:T
16T
13T
01T
1.T
0*T
0)T
0%T
1$T
0#T
1~S
1}S
1|S
1zS
1xS
0'B
0#B
0"B
0~A
0zA
0vA
0sA
0rA
0oA
0nA
0kA
0CU
1AU
0@U
1>U
06U
15U
13U
02U
11U
10U
0,U
0)U
0'U
0~T
0}T
1|T
1#E
0~D
1}D
0|D
0{D
0zD
1yD
0wD
1uD
1tD
0rD
0pD
1oD
1mD
1gD
1fD
1cD
1bD
1`D
1^D
0iU
0hU
0gU
1eU
1dU
1cU
1aU
1[U
1ZU
1YU
0XU
0UU
1SU
0QU
1OU
0MU
1HU
1GU
0oE
0nE
0mE
1lE
0fE
0cE
0_E
0\E
0XE
1UE
0GH
1EH
1DH
0CH
0BH
0AH
1@H
19H
16H
05H
13H
11H
1.H
0%H
0$H
1"H
1}G
0zG
0xG
0wG
0tG
0sG
0rG
0pG
1xH
1uH
0pH
1oH
1lH
0hH
1cH
1_H
0^H
1\H
0YH
0UH
18K
07K
03K
01K
0-K
0,K
0)K
0'K
0&K
0%K
1$K
0"K
0!K
0~J
1{J
0uJ
0sJ
0rJ
1qJ
1jK
1iK
0fK
1eK
1cK
1`K
1^K
1\K
1YK
1XK
1UK
0TK
1SK
1RK
1OK
1NK
1KK
0IK
1HK
0GK
1$W
1}V
0{V
1zV
1vV
0sV
1rV
1nV
1mV
0lV
1kV
0iV
0hV
1gV
0fV
1dV
1`V
1]V
0[V
0RV
1PV
1OV
1GQ
1BQ
1?Q
0;Q
15Q
04Q
0-Q
0)Q
0'Q
1&Q
1}P
0{P
0zP
0xP
1wP
1sP
1rP
1RW
0JW
1GW
1DW
1BW
0=W
1<W
0:W
08W
16W
15W
12W
01W
00W
0-W
1,W
1)W
1(W
0]O
1\O
1XO
1VO
1KO
0JO
1IO
0FO
1dP
1_P
1\P
0XP
1RP
0QP
0JP
0FP
0DP
1CP
1<P
0:P
09P
07P
16P
12P
11P
1FX
1AX
0?X
1>X
1:X
07X
16X
04X
02X
11X
10X
1/X
1-X
0+X
1*X
1)X
0(X
1&X
1!X
0|W
1zW
0xW
0vW
0uW
1tW
0pW
0mW
1lW
1iW
1hW
0GQ
0BQ
0?Q
18Q
07Q
13Q
02Q
01Q
0.Q
1-Q
0,Q
0+Q
1)Q
0~P
0uP
0rP
1TD
0QD
1PD
0OD
0ND
0MD
1LD
0JD
1HD
1GD
0ED
0CD
1BD
1@D
1:D
19D
16D
15D
13D
11D
0=V
1;V
0:V
18V
07V
16V
15V
03V
12V
11V
00V
1-V
1,V
1+V
1*V
0)V
0(V
0'V
1}U
1{U
0yU
0xU
1wU
1vU
1tU
1sU
0#E
1vD
0sD
1pD
1lD
0gD
0`D
0_D
0^D
0a@
1_@
1]@
0Y@
1X@
1U@
0T@
1S@
1P@
1N@
1H@
1F@
0E@
1D@
0vT
0sT
1oT
1mT
0lT
0hT
1fT
1eT
0cT
0aT
1_T
1^T
0\T
0[T
1ZT
1YT
0WT
1VT
0ST
1RT
1OT
1NT
1MT
1KT
1IT
16A
02A
01A
0.A
0,A
0)A
0!A
0y@
0o<
0l<
1k<
1j<
1i<
1h<
0g<
0a<
1`<
1_<
1[<
1Y<
0X<
1T<
1S<
1P<
0ES
0DS
1BS
0@S
0>S
0<S
0;S
09S
07S
06S
15S
13S
12S
0/S
1)S
1'S
1&S
0#S
0"S
1!S
1~R
0}R
0|R
1@=
08=
12=
01=
0-=
1,=
0)=
0#=
0"=
1r<
0j<
1d<
0c<
0_<
1^<
0[<
0U<
0T<
0k=
0j=
1h=
1g=
0f=
0c=
1`=
0]=
0\=
0[=
1W=
0U=
0S=
0Q=
1P=
1O=
0M=
1K=
1I=
1G=
1F=
0E=
0D=
04>
01>
10>
1)>
1(>
0&>
1%>
1~=
1|=
0{=
1x=
0t=
1o=
1d@
0`@
0_@
0\@
0Z@
0W@
0O@
0I@
0hA
0eA
0^A
0]A
1ZA
0YA
0WA
1TA
1QA
1MA
1LA
0KA
1IA
1FA
0AA
1@A
1?A
1=A
1;A
10B
1.B
0+B
1)B
1(B
0%B
1!B
0|A
1zA
0xA
1wA
0tA
1sA
1pA
0TD
1ID
0FD
1CD
1?D
0:D
03D
02D
01D
0QE
1OE
0LE
1HE
0EE
1BE
0@E
1>E
1;E
1:E
04E
11E
10E
1.E
0,E
1+E
1*E
1)E
1xE
0wE
1vE
0tE
0sE
1rE
1qE
0pE
1mE
0jE
0iE
0gE
1`E
1_E
1YE
1XE
0VE
0UE
0dP
0_P
0\P
1UP
0TP
1PP
0OP
0NP
0KP
1JP
0IP
0HP
1FP
0=P
04P
01P
1CO
0BO
1>O
0=O
0<O
1;O
1:O
17O
16O
04O
13O
01O
10O
1.O
0-O
0,O
0*O
0'O
0&O
0%O
1$O
1#O
1"O
1!O
1|N
1yN
0xN
1wN
0vN
0qN
0nN
0jN
1iN
1fN
1eN
1$P
1}O
0vO
0oO
1mO
1lO
1jO
1gO
1fO
0dO
0bO
0[O
1ZO
0WO
0UO
1SO
1PO
1OO
0KO
1BO
1=O
0:O
03O
02O
0.O
1-O
1,O
0)O
1(O
1'O
1&O
0$O
0yN
1pN
0mN
0$P
0}O
1sO
1nO
0mO
0lO
0gO
0fO
1dO
0RO
0NE
1CE
1@E
1=E
09E
14E
1-E
1,E
0+E
0lE
1eE
0`E
0YE
0XE
1dA
1`A
1_A
0\A
0ZA
1WA
0OA
0IA
01B
00B
0(B
1j=
0b=
1\=
1[=
0W=
0V=
1S=
1M=
1L=
0(>
1#>
0~=
0x=
0w=
#82800
b11110100000000000111101011101000 d
b11100010110010100100111011000101 e
0"
1)Y
0(Y
0&Y
1|X
0{X
1yX
0xX
0uX
1tX
0sX
0rX
1pX
0oX
0mX
1u!
0t!
0r!
1j!
0i!
1g!
0f!
0c!
1b!
0a!
0`!
1^!
0]!
0[!
0fX
1dX
0cX
0_X
1^X
1[X
0SX
0RX
0OX
1MX
0LX
1HX
0E!
0C!
0B!
0<!
19!
05!
03!
12!
11!
0.!
1*!
1(!
0%!
0#!
0}
1|
1{
0z
1y
1s
1r
1q
0p
1m
0k
0i
0h
0g
0f
0T!
1r(
0q(
0o(
1g(
0f(
1d(
0c(
0`(
1_(
0^(
0](
1[(
0Z(
0X(
06"
14"
03"
0/"
1."
1+"
0#"
0""
0}!
1{!
0z!
1v!
1zQ
b1 vQ
0tQ
b0 sQ
1qQ
1nQ
b0 jQ
b0 ^Q
1YQ
b1 XQ
b0 LQ
1PQ
b1 OQ
b0 KQ
b111010011010110110001001110101 NQ
b11101001101011011000100111010 QQ
b11101001101011011000100111010 WQ
b11101001101011011000100111010 ZQ
b0 ]Q
b111000101100101001001110110001010 `Q
b0 iQ
b0 lQ
b0 oQ
b111100010110010100100111011000101 rQ
b11101001101011011000100111010 uQ
b0 xQ
1t(
0v(
1w(
1x(
1!)
1$)
0o'
0n'
0m'
0j'
0i'
0g'
0f'
0d'
0a'
0_'
0^'
0\'
0['
0Z'
0X'
0W'
0V'
0S'
0R'
0Q'
1O'
1M'
1L'
1K'
1H'
1D'
1C'
1A'
1@'
1>'
1<'
1;'
18'
16'
15'
14'
0.'
1-'
0*'
1('
1%'
1$'
0#'
0~&
1z&
0y&
1w&
1v&
0u&
1t&
0q&
1o&
1n&
1m&
0k&
0j&
0i&
0f&
0e&
0c&
0b&
0`&
0]&
0[&
0Z&
0X&
0W&
0V&
0T&
0S&
0R&
0O&
0N&
0M&
0L&
0J&
0I&
0H&
0E&
0D&
0B&
0A&
0?&
0<&
0:&
09&
07&
06&
05&
03&
02&
01&
0.&
0-&
0,&
0+&
0*&
0&&
0%&
0"&
0}%
0{%
0z%
0x%
0u%
0q%
0m%
0l%
1$%
0#%
0!%
1w$
0v$
1t$
0s$
0p$
1o$
0n$
0m$
1k$
0j$
0h$
0b$
0^$
0]$
0Z$
0W$
0U$
0T$
0R$
0O$
0K$
0G$
0F$
0A$
1>$
1=$
0;$
19$
08$
14$
03$
11$
00$
1/$
1,$
1'$
1&$
0$$
1}#
0|#
1y#
0w#
0t#
0s#
1r#
1o#
0k#
1j#
0h#
0g#
1f#
0e#
1b#
0`#
0_#
0^#
0<#
1;#
19#
01#
10#
0.#
1-#
1*#
0)#
1(#
1'#
0%#
1$#
1"#
1y"
0x"
0v"
1u"
1t"
0r"
0o"
0m"
1l"
1k"
0j"
1i"
0g"
1f"
0e"
0a"
0_"
1^"
1]"
0["
0Z"
0Y"
0X"
0W"
0S"
0R"
0O"
0L"
0J"
0I"
0G"
0D"
0@"
0<"
0;"
16(
04(
1<(
0@(
0H(
0N(
1P(
0m)
0l)
0h)
0g)
0d)
0a)
0_)
0^)
0\)
0Y)
0U)
0Q)
0P)
1/,
0-,
1,,
1*,
0",
1!,
0}+
1|+
1y+
0x+
1w+
1v+
0t+
1s+
1q+
1-/
0+/
1(/
1'/
0%/
1#/
0"/
1|.
0{.
1y.
0x.
1w.
1t.
1o.
1n.
0l.
0Q/
0M/
0L/
0I/
0F/
0D/
0C/
0A/
0>/
0:/
06/
05/
0y/
1v/
0u/
0s/
1k/
0j/
1h/
0g/
0d/
1c/
0b/
0a/
1_/
0^/
0\/
0u2
0q2
0p2
0m2
0j2
0h2
0g2
0e2
0b2
0^2
0Z2
0Y2
0%8
1"8
1~7
1}7
1|7
1y7
1u7
1t7
1r7
1q7
1o7
1m7
1l7
1i7
1g7
1f7
1e7
03*
11*
00*
0.*
1-*
1,*
0**
0'*
0%*
1$*
1#*
0"*
1!*
0})
1|)
0{)
0w)
0u)
1t)
1s)
0q)
0p)
0o)
1n)
1x,
0w,
1t,
0r,
0o,
0n,
1m,
1j,
0f,
1e,
0c,
0b,
1a,
0`,
1],
0[,
0Z,
0Y,
1X,
0)5
0&5
0%5
0$5
0!5
0~4
0|4
0{4
0y4
0v4
0t4
0s4
0q4
0p4
0o4
0m4
0l4
0k4
0h4
0g4
0f4
0e4
1d4
0L5
0K5
0J5
0G5
0F5
0D5
0C5
0A5
0>5
0<5
0;5
095
085
075
055
045
035
005
0/5
0.5
0-5
1,5
0r5
1q5
0n5
1l5
1i5
1h5
0g5
0d5
1`5
0_5
1]5
1\5
0[5
1Z5
0W5
1U5
1T5
1S5
0R5
1I8
0E8
0D8
0C8
0@8
0?8
0=8
0<8
0:8
078
058
048
028
018
008
0.8
0-8
0,8
0)8
0(8
0'8
1&8
057
027
017
1/7
0,7
0+7
0*7
1)7
0#7
1!7
1|6
0y6
0x6
1w6
0s6
0q6
1m6
0l6
0X7
0W7
0V7
0R7
0Q7
0O7
0J7
0I7
0H7
0G7
0F7
0E7
0C7
0A7
0?7
0<7
0;7
187
0':
1%:
1$:
1":
0}9
0{9
0z9
1y9
0s9
0l9
0j9
0i9
0f9
1c9
1b9
1a9
1`9
1C:
0A:
1;:
11:
0+:
0*:
0):
014
0-4
0,4
0)4
0&4
0$4
0#4
0!4
0|3
0x3
0t3
0s3
191
171
141
131
021
011
101
0.1
0-1
1)1
0(1
0'1
1$1
1#1
0~0
0}0
0z0
0y0
0x0
1w0
0v0
0_1
0]1
1Z1
0Y1
0X1
0Q1
1O1
0N1
0K1
1G1
0F1
1D1
1C1
0B1
0A1
1;.
19.
18.
16.
04.
03.
10.
0-.
0).
1'.
0%.
1$.
1|-
0{-
0z-
1w-
0u-
1t-
0s-
1r-
0a.
1\.
0V.
1U.
0S.
1Q.
1M.
0J.
1I.
0F.
1E.
0>.
0@+
1?+
0>+
1:+
11+
1/+
1,+
0++
1)+
0'+
1#+
0!+
0~*
0}*
0|*
0e+
0`+
0\+
0Y+
0W+
0T+
0Q+
0M+
0I+
1B+
#84600
1"
1T!
b11101001101011011000100111010100 N:
b100000000000000000000000000000000000 O:
b1010111100111001101110101000101001101101 P:
b1000100010001000100010010000000 Q:
b101100100010001111100011010011001101101 R:
b10000001100100000001100100000010000000 S:
b1010100000000000000000000000000000000000 T:
b101000010110010100100111011000101000000 V:
b10100000000000000000000000000000000000 W:
b11110100100001100000111001000011101100 X:
b1010100010101000100010000000000 Y:
b111111110110010000011110001100010111100 "F
b10000000001001001010100010010001000000000 #F
b1010110000010001011100101111100000001110110000 $F
b1001000100100001000000010010100000000000 %F
b11101111110010011011111110110000110000011001 &F
b10001101100100000001000110001010000000 'F
b100000010110001000001110011100111110010110001110 xK
b1001010010101010100011001000101001000000 yK
b1101110001000001110100000010001011000010000100100000000 zK
b100101110011011011101010100101000110000000000000 {K
b1101100101000010100001001010111100111000110010000011010101110011 HQ
b10000011001001010101001000010001010001000010000000000000000 IQ
b101011110011101100100100010110100111000010100010010001000 P!
b1111010001100010011010010101110000010110100101010000110010111100 Q!
b1101111010011111001011100101100001110111000111101111101000001110 R!
b1110000101110100110110011101000001001101000010100011010101110011 S!
b11110100000000000111101011101000 H!
b1111001001100000110100111110010 J!
b10001001001100101101011000010010 L!
b1110010101011111111011111100101 N!
b11100010110010100100111011000101 I!
b11100111011101101001011011001110 K!
b1000111111011001101101110001111 M!
b10111011110100100111001001110111 O!
0hY
1eY
1dY
1bY
0`Y
1_Y
0]Y
0\Y
0[Y
0ZY
1YY
0XY
0VY
1RY
0QY
0LY
0KY
1GY
1AY
0@Y
0?Y
1;Y
09Y
07Y
06Y
05Y
14Y
13Y
02Y
00Y
0.Y
1,Y
1c
1^
0\
1[
1W
1V
0U
0T
0Q
1P
0N
0M
0L
1K
0J
1H
1E
0D
0C
0A
0@
1?
0>
1=
1<
09
17
06
15
14
02
00
1.
0,
1+
0)
1&
1%
1$
1JN
1IN
0FN
1EN
1CN
1@N
1>N
1<N
19N
18N
15N
04N
13N
12N
1/N
1.N
1+N
0)N
1(N
0'N
1nM
0mM
0iM
0gM
0cM
0bM
0_M
0]M
0\M
0[M
1ZM
0XM
0WM
0VM
1SM
0MM
0KM
0JM
1IM
18M
15M
00M
1/M
1,M
0(M
1#M
1}L
0|L
1zL
0wL
0sL
0]L
1[L
1ZL
0YL
0XL
0WL
1VL
1OL
1LL
0KL
1IL
1GL
1DL
0;L
0:L
18L
15L
02L
00L
0/L
0,L
0+L
0*L
0(L
1TJ
0SJ
1RJ
0PJ
0OJ
1NJ
1MJ
0LJ
0KJ
0JJ
0FJ
0EJ
0CJ
0BJ
1AJ
0?J
08J
04J
02J
0#J
1!J
0~I
0|I
1xI
0uI
1sI
1rI
1nI
1mI
1kI
1jI
0iI
1aI
1`I
1^I
1]I
1ZI
1YI
0OI
1LI
0II
1GI
0EI
0CI
0AI
0@I
1?I
0>I
0<I
08I
17I
06I
04I
02I
10I
0/I
0.I
0+I
0fG
0cG
1bG
1^G
1]G
0\G
0[G
0ZG
0WG
1RG
1OG
0MG
1KG
1JG
0IG
1DG
0?G
1>G
1=G
1;G
19G
01G
0.G
1-G
0(G
1&G
1~F
0zF
1yF
0xF
0qF
0nF
1lF
0]F
1ZF
1YF
0XF
0UF
0TF
1RF
0OF
0HF
0GF
0CF
1BF
1AF
1>F
1=F
1;F
19F
18F
07F
06F
1zC
0xC
1rC
1hC
0bC
0aC
0`C
0YC
1WC
1VC
1TC
0QC
0OC
0NC
1MC
0GC
0@C
0>C
0=C
0:C
17C
16C
15C
14C
0-C
0,C
0+C
0'C
0&C
0$C
0}B
0|B
0{B
0zB
0yB
0xB
0vB
0tB
0rB
0oB
0nB
1kB
0eB
0bB
0aB
1_B
0\B
0[B
0ZB
1YB
0SB
1QB
1NB
0KB
0JB
1IB
0EB
0CB
1?B
0>B
0\?
0X?
0W?
0T?
0Q?
0O?
0N?
0L?
0I?
0E?
0A?
0@?
06?
04?
11?
00?
0/?
0(?
1&?
0%?
0"?
1|>
0{>
1y>
1x>
0w>
0v>
1h>
1f>
1c>
1b>
0a>
0`>
1_>
0]>
0\>
1X>
0W>
0V>
1S>
1R>
0O>
0N>
0K>
0J>
0I>
1H>
0G>
0D<
1?<
09<
18<
06<
14<
10<
0-<
1,<
0)<
1(<
0!<
1z;
1x;
1w;
1u;
0s;
0r;
1o;
0l;
0h;
1f;
0d;
1c;
1];
0\;
0[;
1X;
0V;
1U;
0T;
1S;
0P;
0K;
0G;
0D;
0B;
0?;
0<;
08;
04;
1-;
0%;
1$;
0#;
1}:
1t:
1r:
1o:
0n:
1l:
0j:
1f:
0d:
0c:
0b:
0a:
1LR
0KR
1HR
1GR
0DR
0AR
1?R
1>R
08R
16R
05R
04R
11R
10R
0.R
0-R
0,R
0+R
1*R
0@=
1?=
1==
1:=
07=
14=
11=
1+=
1)=
1(=
1#=
1"=
0!=
0~<
1wR
1uR
1rR
0pR
0lR
0hR
1fR
0eR
0dR
1cR
0aR
0]R
0\R
1ZR
1UR
0SR
1RR
1PR
1/>
0)>
1$>
1v=
0o=
1vS
1tS
1sS
1pS
0oS
1lS
0kS
0jS
1fS
1dS
1cS
1bS
1aS
1`S
1_S
0]S
0\S
1[S
1ZS
0YS
0;T
07T
06T
03T
00T
0.T
0-T
0+T
0(T
0$T
0~S
0}S
19A
17A
13A
0-A
1)A
0(A
0'A
1$A
1#A
0~@
0}@
0x@
0v@
0t@
0EU
0BU
0AU
0>U
1=U
0<U
0;U
0:U
18U
16U
03U
00U
0/U
0-U
1,U
0+U
1)U
1(U
1&U
0%U
0"U
0|T
0!E
1|D
1zD
0uD
0tD
1sD
0mD
0jD
1iD
0cD
1_D
0kU
1iU
1hU
1fU
0cU
0aU
1_U
0^U
0YU
1XU
0RU
1PU
0OU
0NU
1LU
1IU
1nE
1fE
1\E
0FH
1CH
1BH
0?H
1<H
07H
15H
14H
03H
01H
10H
1+H
1(H
1'H
0!H
0}G
1|G
1{G
0vG
1uG
1tG
1rG
1pG
0xH
0uH
0sH
1rH
0oH
1nH
1mH
0lH
0kH
0gH
0cH
1bH
1[H
1XH
0WH
08K
05K
13K
12K
11K
1-K
0+K
1'K
1&K
1%K
1#K
1!K
1}J
1|J
0yJ
0xJ
0wJ
1uJ
1rJ
0qJ
1pJ
1oJ
1nJ
0mJ
0kJ
1jJ
1lK
0jK
0iK
0eK
0cK
1bK
0`K
0^K
0\K
0ZK
0XK
1WK
0VK
0UK
0RK
1QK
1PK
0OK
0NK
0KK
1JK
0HK
1FK
0$W
1"W
1!W
0~V
0}V
0|V
0xV
1tV
1sV
0rV
1qV
0pV
1oV
0nV
1lV
0kV
1iV
1fV
1bV
1aV
0`V
0]V
1\V
0ZV
0XV
0WV
0UV
0TV
0QV
0PV
0OV
0MV
1EQ
1DQ
1@Q
19Q
16Q
05Q
11Q
0/Q
1.Q
0%Q
0$Q
1"Q
0}P
0sP
0pP
1SW
0RW
0NW
1MW
0IW
0GW
0FW
0DW
0CW
0BW
0@W
1=W
07W
06W
05W
11W
10W
0/W
0,W
1+W
1*W
1kO
0hO
1eO
1`O
1[O
1WO
0VO
1UO
1TO
1QO
1MO
1JO
0IO
1bP
1aP
1]P
1VP
1SP
0RP
1NP
0LP
1KP
0BP
0AP
1?P
0<P
02P
0/P
0FX
1DX
1CX
0BX
0AX
0@X
0<X
18X
17X
06X
13X
12X
0-X
1+X
0*X
0)X
1(X
0"X
0!X
1~W
1}W
1|W
0zW
1yW
1uW
0sW
1rW
1pW
0lW
1kW
1jW
0EQ
0DQ
1=Q
09Q
08Q
17Q
01Q
0!Q
1}P
0wP
0RD
1OD
1MD
0HD
0GD
1FD
0@D
0=D
1<D
06D
12D
0?V
0<V
0;V
19V
08V
05V
02V
01V
10V
1/V
0,V
0*V
1)V
0%V
1#V
1"V
0}U
1|U
0{U
1xU
0vU
1uU
0|D
0zD
0vD
0sD
0pD
0oD
0lD
0iD
0fD
0bD
1g@
1e@
1a@
0[@
1W@
0V@
0U@
1R@
1Q@
0N@
0M@
0H@
0F@
0D@
1vT
1tT
1sT
1pT
0oT
1lT
0kT
0eT
1dT
1cT
1aT
1`T
1[T
0YT
1WT
1ST
0OT
0NT
09A
07A
06A
03A
0/A
0)A
0%A
0$A
0#A
0"A
0{@
0r<
1q<
1o<
1l<
0i<
1f<
1c<
1]<
1[<
1Z<
1U<
1T<
0S<
0R<
0CS
0BS
1@S
0=S
1<S
17S
16S
05S
03S
02S
11S
0-S
1,S
0*S
0(S
0'S
0&S
1%S
1$S
1#S
0~R
1}R
1{R
0;=
04=
02=
01=
0+=
0)=
0(=
0'=
0}<
0|<
1{<
0m<
0f<
0d<
0c<
0]<
0[<
0Z<
0Y<
0Q<
0P<
1O<
0j=
0h=
0g=
1f=
1d=
1c=
1b=
0a=
1^=
1]=
0\=
0Y=
1X=
1W=
1U=
0P=
1N=
0I=
0F=
1E=
1C=
14>
00>
0/>
1)>
1(>
0%>
0$>
1~=
1}=
0y=
0v=
1t=
0g@
0e@
0d@
0a@
0]@
0W@
0S@
0R@
0Q@
0P@
0K@
1hA
1gA
1fA
1bA
1^A
1]A
1[A
0SA
0QA
0NA
1KA
1IA
1HA
0FA
1EA
1DA
1AA
0@A
16B
0.B
0,B
1$B
1#B
1"B
0zA
0wA
0sA
0pA
0OD
0MD
0ID
0FD
0CD
0BD
0?D
0<D
09D
05D
0SE
0PE
0OE
1ME
1GE
1FE
1EE
1DE
0CE
0BE
1AE
0>E
0=E
0:E
19E
13E
12E
01E
00E
0.E
1+E
0xE
0rE
0qE
1oE
0mE
1jE
1iE
0eE
0_E
0^E
0bP
0aP
1ZP
0VP
0UP
1TP
0NP
0>P
1<P
06P
0CO
1AO
0>O
0=O
0;O
09O
15O
13O
11O
1/O
0,O
1)O
0(O
0'O
0&O
1%O
0~N
0|N
0zN
1yN
1xN
0wN
1vN
0rN
0pN
1oN
1nN
1mN
0kN
0iN
1hN
1gN
1"P
1{O
1tO
0sO
1lO
0jO
1hO
1gO
0eO
0_O
1^O
1]O
0[O
0ZO
0XO
0QO
0PO
0OO
0JO
1@O
0?O
18O
14O
03O
12O
1,O
1zN
0xN
1rN
0"P
0tO
0lO
0\O
1ZO
0TO
0IE
0GE
1CE
0@E
1=E
0<E
09E
16E
03E
0/E
0oE
0iE
0bE
0gA
1eA
0dA
0aA
0]A
0WA
1SA
1RA
1QA
1PA
0KA
06B
0$B
0#B
0"B
0!B
0e=
0^=
1\=
0[=
0U=
0S=
1R=
1Q=
1I=
0H=
0G=
0)>
0}=
0|=
0t=
1r=
#86400
b101110010110000100100101011100 d
b11011110100011100010100010111101 e
0"
1&Y
1%Y
1$Y
0#Y
0~X
0}X
1zX
0yX
1uX
0qX
1mX
1lX
1kX
0jX
1r!
1q!
1p!
0o!
0l!
0k!
1h!
0g!
1c!
0_!
1[!
1Z!
1Y!
0X!
1eX
1cX
0bX
0`X
1_X
0^X
0[X
0ZX
1TX
1SX
1QX
1NX
1LX
0KX
0IX
0HX
1E!
1B!
1A!
0=!
1<!
09!
18!
07!
15!
14!
01!
1/!
1.!
0-!
1,!
1)!
0(!
1&!
1#!
0!!
1~
0{
0y
0x
0w
0s
0r
1p
1n
1j
1i
1h
1g
1f
0T!
1o(
1n(
1m(
0l(
0i(
0h(
1e(
0d(
1`(
0\(
1X(
1W(
1V(
0U(
15"
13"
02"
00"
1/"
0."
0+"
0*"
1$"
1#"
1!"
1|!
1z!
0y!
0w!
0v!
0zQ
b1 pQ
1tQ
0nQ
b1 gQ
0kQ
0_Q
0YQ
b0 XQ
0VQ
0SQ
b0 RQ
b100001011100011101011101000010 NQ
b110111101000111000101000101111010 QQ
b111011110100011100010100010111101 TQ
b111011110100011100010100010111101 WQ
b1000010111000111010111010000101 ZQ
b111011110100011100010100010111101 ]Q
b111011110100011100010100010111101 `Q
b1000010111000111010111010000101 fQ
b110111101000111000101000101111010 iQ
b111011110100011100010100010111101 lQ
b1000010111000111010111010000101 oQ
b0 rQ
b100001011100011101011101000010 uQ
b111011110100011100010100010111101 xQ
0t(
1v(
0x(
0y(
0}(
0!)
0")
0#)
1q'
1o'
1n'
1m'
1l'
1j'
1f'
1d'
1`'
1_'
1^'
1Z'
1X'
1W'
1V'
1U'
1S'
1R'
1Q'
0M'
0L'
0K'
1J'
1G'
1F'
0C'
1B'
0>'
1:'
06'
05'
04'
13'
0/'
0-'
0)'
0('
0&'
0%'
0$'
0!'
0|&
0z&
0w&
0v&
0t&
0p&
0o&
0n&
0m&
1l&
1j&
1e&
1c&
1b&
1a&
1_&
1]&
1\&
1[&
1W&
1V&
1U&
1S&
1N&
1K&
1I&
1H&
1G&
1F&
1D&
1@&
1>&
1:&
19&
18&
14&
12&
11&
10&
1/&
1-&
1,&
1+&
1)&
1'&
1&&
1%&
1$&
1"&
1|%
1z%
1v%
1u%
1t%
1p%
1n%
1m%
1l%
1k%
1i%
1h%
1g%
1e%
1`%
1^%
1]%
1\%
1Z%
1X%
1W%
1V%
1R%
1Q%
1P%
1N%
1I%
1%%
0$%
1#%
1!%
1~$
0{$
0y$
0w$
1v$
0t$
1r$
1p$
0o$
0k$
1j$
1h$
1g$
1b$
1`$
1_$
1^$
1]$
1[$
1W$
1U$
1Q$
1P$
1O$
1K$
1I$
1H$
1G$
1F$
1D$
1C$
1B$
1A$
0@$
1?$
0>$
0=$
0<$
1:$
09$
18$
17$
16$
05$
10$
0/$
0-$
1+$
1*$
0)$
1($
0'$
0&$
0%$
1#$
1~#
0}#
1|#
1w#
0v#
1s#
0r#
0o#
0n#
1m#
1k#
0j#
0i#
1g#
0f#
1e#
1`#
1_#
1^#
1]#
1[#
1Z#
1Y#
1X#
1V#
1R#
1P#
1L#
1K#
1J#
1F#
1D#
1C#
1B#
1A#
1?#
1>#
1=#
16#
0/#
1.#
0-#
0,#
1)#
0'#
1}"
1{"
1z"
0y"
1x"
0w"
0u"
0t"
1q"
1o"
1m"
0l"
1j"
0h"
0f"
1e"
1a"
0`"
0^"
0]"
08(
0<(
1F(
1L(
01*
10*
0/*
0-*
0,*
1)*
1'*
1%*
0$*
1"*
0~)
0|)
1{)
1w)
0v)
0t)
0s)
0-/
1+/
0*/
1)/
0(/
0'/
0&/
1$/
0#/
1"/
1!/
1~.
0}.
1x.
0w.
0u.
1s.
1r.
0q.
1p.
0o.
0n.
0m.
1k.
1w/
0v/
1u/
1s/
1r/
0o/
0m/
0k/
1j/
0h/
1f/
1d/
0c/
0_/
1^/
1\/
1[/
1O2
1M2
1H2
1F2
1E2
1D2
1B2
1@2
1?2
1>2
1:2
192
182
162
112
1M5
1K5
1F5
1D5
1C5
1B5
1@5
1>5
1=5
1<5
185
175
165
145
1/5
0~7
0}7
0|7
1{7
1x7
1w7
0t7
1s7
0o7
1k7
0g7
0f7
0e7
1d7
1',
0~+
1}+
0|+
0{+
1x+
0v+
1n+
1l+
1k+
0j+
0U,
1S,
1Q,
1P,
1O,
1N,
1L,
1H,
1F,
1B,
1A,
1@,
1<,
1:,
19,
18,
17,
15,
14,
13,
02,
1y,
0x,
1w,
1r,
0q,
1n,
0m,
0j,
0i,
1h,
1f,
0e,
0d,
1b,
0a,
1`,
1[,
1Z,
1Y,
0X,
1Q/
1O/
1N/
1M/
1L/
1J/
1F/
1D/
1@/
1?/
1>/
1:/
18/
17/
16/
15/
13/
12/
11/
00/
1w2
1t2
1r2
1q2
1p2
1o2
1m2
1i2
1g2
1c2
1b2
1a2
1]2
1[2
1Z2
1Y2
1X2
1V2
1U2
0T2
1'5
1%5
1$5
1#5
1"5
1~4
1z4
1x4
1t4
1s4
1r4
1n4
1l4
1k4
1j4
1i4
1g4
1f4
1e4
0d4
1u5
0s5
0q5
0m5
0l5
0j5
0i5
0h5
0e5
0b5
0`5
0]5
0\5
0Z5
0V5
0U5
0T5
0S5
1R5
1G8
1E8
1D8
1C8
1B8
1@8
1<8
1:8
168
158
148
108
1.8
1-8
1,8
1+8
1)8
1(8
1'8
0&8
09.
17.
13.
02.
00.
1..
1-.
1+.
0*.
0&.
0$.
1".
1!.
1z-
0y-
0x-
1s-
0r-
1].
1[.
1Z.
1X.
0U.
1R.
0Q.
1N.
1L.
0I.
1F.
1D.
1C.
1B.
1A.
1?.
1#:
0":
1|9
0y9
0u9
0t9
1q9
1p9
1o9
0n9
0m9
1j9
1i9
0e9
0c9
0b9
0a9
0`9
1E:
1B:
1A:
1=:
1<:
09:
16:
15:
01:
1.:
1-:
1+:
1*:
1):
137
117
107
0/7
1.7
0-7
1,7
1*7
0)7
0(7
1'7
0&7
0%7
0!7
0|6
0z6
1y6
0v6
1u6
0t6
1s6
1r6
0o6
1n6
0m6
1l6
1Y7
1W7
1P7
1N7
1J7
1I7
1H7
1D7
1B7
1@7
1;7
0:7
087
114
104
1.4
1-4
1+4
1*4
1(4
1&4
1%4
1$4
1"4
1}3
1z3
1x3
1w3
1u3
1t3
0r3
0p3
1o3
0n3
1[4
1T4
1Q4
1K4
1F4
1E4
1=4
1<4
1:4
091
071
061
041
031
121
1.1
1-1
0,1
0*1
0)1
1(1
1'1
0%1
0!1
0{0
1y0
1v0
0t0
0s0
1r0
1_1
1]1
1[1
0Z1
1Y1
1X1
1V1
1T1
0S1
1R1
0O1
1N1
1J1
1I1
1H1
0G1
1F1
0C1
1B1
1A1
1?1
1>1
1=1
0<1
0?+
1>+
0=+
0;+
0:+
17+
15+
13+
02+
10+
0.+
0,+
1++
1'+
0&+
0$+
0#+
#88200
1"
1T!
b10000101110001110101110100001000 N:
b110110010111111000110011110000101111001 P:
b1011111100000111000100000111111000000 Q:
b110001101000000111001100001111010000000 R:
b1110110101011100010101010101101010100 S:
b100001101101001001011101011011011000000 T:
b10110000000110000100000100100000010000 U:
b1010001101010100000000100100101010110100 V:
b10000101010001110001010000001010000 W:
b111000011100001000001011011100 X:
b1110111000101110001110101110100000000 Y:
b101000111111101100001101011001011101001000 "F
b10000000000011010000100010000000100000 #F
b1010101001100111011001111111000010011101101101 $F
b10000000000000000 %F
b11111100001010111001010101011110100001000000 &F
b10100001000010001000100000001000000000 'F
b101011000001100010001110011110101011101110110010111100 xK
b101110010110010000000110001000000000000 yK
b1110101110100100000111010111111010010011110000000000000 zK
b10001001001101000101000000001000000000100000000000 {K
b1101111000011100100010011000011101000100110111101111100000001110 HQ
b1000001010100100110100010011001001000000000000100000000 IQ
b1111100111110010000000101001101001111011101011001000100011101100 P!
b101011110011101100100100010110100111000010100010010001000 Q!
b1111010001100010011010010101110000010110100101010000110010111100 R!
b1101111010011111001011100101100001110111000111101111101000001110 S!
b101110010110000100100101011100 H!
b11110100000000000111101011101000 J!
b1111001001100000110100111110010 L!
b10001001001100101101011000010010 N!
b11011110100011100010100010111101 I!
b11100010110010100100111011000101 K!
b11100111011101101001011011001110 M!
b1000111111011001101101110001111 O!
0gY
0eY
0dY
0^Y
1[Y
0WY
0UY
1TY
1SY
0PY
1LY
1JY
0GY
0EY
0AY
1@Y
1?Y
0>Y
1=Y
17Y
16Y
15Y
04Y
11Y
0/Y
0-Y
0,Y
0+Y
0*Y
0c
1a
1`
0_
0^
0]
0[
1Z
0Y
1X
1U
1T
1Q
1O
1J
0H
1G
1F
1@
0<
0;
1:
19
07
16
05
04
13
12
10
0.
0-
1,
0+
1*
1)
1(
1'
0&
1LN
0JN
0IN
0EN
0CN
1BN
0@N
0>N
0<N
0:N
08N
17N
06N
05N
02N
11N
10N
0/N
0.N
0+N
1*N
0(N
1&N
0nM
0kM
1iM
1hM
1gM
1cM
0aM
1]M
1\M
1[M
1YM
1WM
1UM
1TM
0QM
0PM
0OM
1MM
1JM
0IM
1HM
1GM
1FM
0EM
0CM
1BM
08M
05M
03M
12M
0/M
1.M
1-M
0,M
0+M
0'M
0#M
1"M
1yL
1vL
0uL
0\L
1YL
1XL
0UL
1RL
0ML
1KL
1JL
0IL
0GL
1FL
1AL
1>L
1=L
07L
05L
14L
13L
0.L
1-L
1,L
1*L
1(L
0TJ
0NJ
0MJ
1JJ
0IJ
1FJ
1BJ
0AJ
0>J
0;J
0:J
18J
0%J
0"J
0!J
1}I
0yI
1vI
1uI
1tI
0rI
1qI
0pI
0nI
0lI
0jI
1fI
1bI
0aI
0`I
0_I
0^I
1[I
0LI
0JI
0?I
0:I
07I
03I
00I
1fG
1dG
1cG
0bG
1`G
0_G
1\G
1YG
0UG
1PG
1NG
0LG
1GG
1FG
0DG
1CG
1BG
1?G
0>G
11G
0-G
0&G
1%G
0"G
1{F
0yF
0vF
1oF
0lF
0\F
0ZF
0YF
1XF
0WF
1VF
1UF
1TF
0SF
1OF
0MF
0KF
1JF
1IF
0EF
1DF
1CF
0BF
1@F
0:F
09F
08F
17F
15F
1|C
1yC
1xC
1tC
1sC
0pC
1mC
1lC
0hC
1eC
1dC
1bC
1aC
1`C
1UC
0TC
1PC
0MC
0IC
0HC
1EC
1DC
1CC
0BC
0AC
1>C
1=C
09C
07C
06C
05C
04C
1.C
1,C
1%C
1#C
1}B
1|B
1{B
1wB
1uB
1sB
1nB
0mB
0kB
1cB
1aB
1`B
0_B
1^B
0]B
1\B
1ZB
0YB
0XB
1WB
0VB
0UB
0QB
0NB
0LB
1KB
0HB
1GB
0FB
1EB
1DB
0AB
1@B
0?B
1>B
1.@
1'@
1$@
1|?
1w?
1v?
1n?
1m?
1k?
1\?
1[?
1Y?
1X?
1V?
1U?
1S?
1Q?
1P?
1O?
1M?
1J?
1G?
1E?
1D?
1B?
1A?
0??
0=?
1<?
0;?
16?
14?
12?
01?
10?
1/?
1-?
1+?
0*?
1)?
0&?
1%?
1!?
1~>
1}>
0|>
1{>
0x>
1w>
1v>
1t>
1s>
1r>
0q>
0h>
0f>
0e>
0c>
0b>
1a>
1]>
1\>
0[>
0Y>
0X>
1W>
1V>
0T>
0P>
0L>
1J>
1G>
0E>
0D>
1C>
1@<
1><
1=<
1;<
08<
15<
04<
11<
1/<
0,<
1)<
1'<
1&<
1%<
1$<
1"<
0x;
1v;
1r;
0q;
0o;
1m;
1l;
1j;
0i;
0e;
0c;
1a;
1`;
1[;
0Z;
0Y;
1T;
0S;
0$;
1#;
0";
0~:
0}:
1z:
1x:
1v:
0u:
1s:
0q:
0o:
1n:
1j:
0i:
0g:
0f:
0LR
1KR
0JR
0HR
0GR
1DR
1BR
1@R
0?R
1=R
0;R
09R
18R
14R
03R
01R
00R
1>=
0==
1;=
17=
06=
15=
13=
12=
11=
10=
1/=
0.=
1+=
0*=
1'=
1&=
0uR
1sR
1pR
0oR
1mR
1lR
1kR
1jR
1iR
1hR
1gR
0fR
1eR
1dR
0bR
1aR
1`R
0_R
1^R
1]R
1\R
1YR
0XR
0UR
0TR
0RR
1QR
0PR
10>
1.>
1->
1+>
0(>
1%>
1w=
1s=
0vS
0tS
0pS
0nS
0mS
0lS
1kS
0iS
1hS
1eS
0dS
0cS
1]S
1\S
0[S
0XS
0WS
0VS
1PS
12A
1.A
1-A
1,A
0*A
1)A
1(A
1'A
1&A
1$A
1"A
1!A
1|@
1y@
1v@
1t@
1s@
1r@
1<T
1;T
1:T
18T
17T
14T
10T
1/T
1.T
1)T
1'T
1$T
1#T
1!T
1~S
1{S
0zS
0xS
1.B
1vA
1mA
1kA
1CU
1AU
0?U
0=U
1<U
1:U
09U
08U
06U
10U
1/U
0.U
0,U
0)U
0(U
0&U
1%U
1$U
1"U
1~T
1|T
1%E
1#E
1"E
1~D
1|D
1zD
1wD
1vD
0nD
1kD
1iD
0hD
1gD
1eD
1dD
0aD
1`D
0_D
1^D
1gU
0fU
1^U
0[U
1YU
1WU
1UU
1TU
1RU
0PU
1OU
1NU
1JU
0IU
1lE
1hE
1gE
0\E
1XE
0EH
0CH
0BH
0@H
1>H
0=H
1;H
09H
04H
13H
02H
0,H
0(H
0'H
1%H
1#H
0"H
1}G
0{G
1zG
1yG
1vG
0uG
1xH
1vH
1tH
0rH
1pH
0mH
1lH
1iH
0eH
1dH
1cH
0bH
1`H
1^H
0\H
0ZH
1WH
03K
02K
01K
1/K
0-K
1+K
0$K
0#K
0}J
0|J
1yJ
1xJ
1wJ
1vJ
0uJ
0pJ
0nJ
1kJ
0lK
0bK
1ZK
0YK
0WK
1VK
0SK
0QK
0PK
0JK
0#W
1~V
1}V
1{V
0zV
1xV
1wV
0vV
0uV
0qV
0lV
1kV
0jV
1eV
1cV
0bV
1^V
0\V
1[V
1YV
1XV
0SV
1RV
1QV
1OV
1MV
1CQ
1BQ
1<Q
07Q
06Q
15Q
03Q
11Q
10Q
1/Q
1+Q
0)Q
1(Q
1$Q
1!Q
0}P
1|P
1{P
0vP
1uP
1tP
1rP
1pP
0SW
0PW
1OW
1NW
0EW
1CW
1BW
1@W
1?W
1>W
0=W
0<W
0;W
18W
16W
13W
01W
1/W
1,W
0*W
0)W
0(W
1'W
0kO
0gO
0`O
0^O
1YO
0WO
1RO
0MO
1LO
1`P
1_P
1YP
0TP
0SP
1RP
0PP
1NP
1MP
1LP
1HP
0FP
1EP
1AP
1>P
0<P
1;P
1:P
05P
14P
13P
11P
1/P
0EX
1BX
1AX
1?X
0>X
1<X
1;X
0:X
09X
02X
01X
0/X
1.X
1)X
0&X
0%X
1$X
1!X
0|W
1zW
1xW
1vW
0uW
0tW
1lW
0jW
0iW
0hW
1gW
0CQ
0BQ
0@Q
0=Q
0<Q
1:Q
16Q
01Q
0/Q
1'Q
1#Q
0!Q
0|P
0uP
0tP
0rP
1VD
1TD
1SD
1QD
1OD
1MD
1JD
1ID
0AD
1>D
1<D
0;D
1:D
18D
17D
04D
13D
02D
11D
1=V
1;V
09V
17V
06V
15V
13V
12V
00V
1,V
1*V
1(V
1'V
1&V
1%V
1}U
1{U
0xU
0uU
0%E
0#E
0}D
0zD
0yD
0xD
0vD
1pD
0eD
1bD
0`D
0^D
1`@
1\@
1[@
1Z@
0X@
1W@
1V@
1U@
1T@
1R@
1P@
1O@
1L@
1I@
1F@
1D@
1C@
1B@
0vT
0tT
0pT
0nT
0mT
0lT
1jT
1hT
1gT
0fT
1eT
0dT
0_T
0^T
1\T
0[T
0WT
0ST
0RT
1OT
1LT
0KT
0IT
10A
1/A
0.A
0,A
0(A
0&A
1~@
0|@
1w@
1p<
0o<
1m<
1i<
0h<
1g<
1e<
1d<
1c<
1b<
1a<
0`<
1]<
0\<
1Y<
1X<
1DS
1CS
1?S
1=S
19S
06S
04S
12S
00S
1/S
0.S
1-S
1*S
1(S
1&S
0%S
1"S
0!S
0}R
1|R
0{R
0?=
0>=
0;=
0:=
05=
03=
02=
0,=
0&=
0$=
0#=
0q<
0p<
0m<
0l<
0g<
0e<
0d<
0^<
0X<
0V<
0U<
1j=
0i=
1h=
1g=
0c=
1a=
0`=
0]=
1[=
1Y=
1V=
1S=
0Q=
0N=
0L=
0K=
1H=
1G=
0E=
1D=
0C=
16>
04>
12>
1*>
0%>
0#>
1">
0~=
1|=
1{=
1y=
1v=
0s=
1p=
1^@
1]@
0\@
0Z@
0V@
0T@
1N@
0L@
1G@
0hA
0fA
0bA
0_A
0^A
0[A
1YA
0UA
0TA
0RA
0QA
1OA
1NA
0MA
0LA
1FA
0EA
1CA
1BA
0AA
1>A
0=A
0;A
1-B
1,B
1+B
0)B
1(B
1'B
1&B
1%B
1#B
1|A
1{A
1pA
0mA
0VD
0TD
0PD
0MD
0LD
0KD
0ID
1CD
08D
15D
03D
01D
1QE
1PE
1OE
1NE
1JE
0FE
0CE
1@E
1>E
1<E
1:E
19E
08E
06E
15E
04E
13E
02E
0-E
0,E
1wE
0vE
1uE
1sE
1rE
1pE
1oE
0lE
0jE
0hE
0gE
0fE
1dE
1bE
0aE
1`E
1^E
1]E
1YE
0`P
0_P
0]P
0ZP
0YP
1WP
1SP
0NP
0LP
1DP
1@P
0>P
0;P
04P
03P
01P
0BO
1?O
1=O
1<O
1;O
19O
08O
06O
02O
01O
00O
0/O
1*O
1$O
0"O
0!O
1}N
1|N
0zN
0yN
1xN
0vN
1uN
1sN
0rN
1pN
0oN
0mN
1kN
1iN
0gN
0fN
0eN
1dN
1~O
0{O
1xO
1pO
1kO
1fO
0dO
1aO
1\O
1[O
0ZO
1XO
0UO
1QO
1OO
1HO
1>O
0=O
0;O
18O
07O
05O
11O
0,O
0*O
1"O
0|N
1zN
1wN
0pN
1oN
1mN
0~O
0xO
1uO
1^O
0\O
0YO
0QO
0OO
0PE
0NE
0JE
1GE
1FE
0EE
1CE
0=E
12E
1/E
1-E
0+E
0sE
0rE
0oE
1iE
0^E
0YE
1^A
1]A
1\A
1ZA
0VA
1TA
0NA
1LA
1GA
0-B
0+B
0%B
1}A
0{A
1i=
0h=
1e=
0d=
1_=
1]=
0\=
0V=
1P=
1N=
0M=
06>
02>
0,>
0*>
0{=
0y=
#90000
b10010110101010110101100000101101 d
b10110010101001110010011001100101 e
0"
0&Y
0%Y
1#Y
0"Y
1~X
1}X
0|X
1wX
0tX
1rX
0mX
0lX
1jX
0iX
0r!
0q!
1o!
0n!
1l!
1k!
0j!
1e!
0b!
1`!
0[!
0Z!
1X!
0W!
1gX
0cX
1bX
0aX
0_X
1[X
1WX
1VX
0SX
1RX
0QX
1PX
0LX
1KX
0JX
1HX
1G!
0E!
0D!
0B!
1?!
1>!
1=!
0<!
1;!
1:!
19!
08!
17!
16!
05!
02!
00!
0/!
0.!
0,!
0)!
1(!
0&!
1%!
0~
1}
0|
1{
1u
0p
1l
1k
0h
0g
0f
0T!
0o(
0n(
1l(
0k(
1i(
1h(
0g(
1b(
0_(
1](
0X(
0W(
1U(
0T(
17"
03"
12"
01"
0/"
1+"
1'"
1&"
0#"
1""
0!"
1~!
0z!
1y!
0x!
1v!
1zQ
b1 yQ
0tQ
0wQ
b0 vQ
1nQ
b1 mQ
1kQ
b1 jQ
b1 dQ
1YQ
1SQ
b1 RQ
0MQ
b110110010101001110010011001100101 KQ
b1001101010110001101100110011010 NQ
b1001101010110001101100110011010 QQ
b110110010101001110010011001100101 TQ
b0 WQ
b10011010101100011011001100110101 ZQ
b101100101010011100100110011001010 ]Q
b110110010101001110010011001100101 `Q
b1001101010110001101100110011010 cQ
b1001101010110001101100110011010 fQ
b1001101010110001101100110011010 iQ
b1001101010110001101100110011010 lQ
b1001101010110001101100110011010 oQ
b101100101010011100100110011001010 rQ
b110110010101001110010011001100101 uQ
b10011010101100011011001100110101 xQ
1t(
0v(
0u(
1x(
1y(
1!)
1#)
0%)
0n'
0j'
1i'
1h'
0f'
1e'
1b'
1a'
0`'
0_'
0^'
1]'
1\'
0W'
0S'
0Q'
1P'
0O'
1N'
1K'
0H'
0D'
1C'
0B'
0A'
1?'
1>'
0<'
0:'
19'
08'
17'
14'
11'
10'
1.'
1,'
1)'
1('
1%'
1$'
1!'
1|&
1{&
1z&
1w&
1u&
1s&
1p&
1o&
1m&
0l&
1k&
0j&
1i&
1h&
1d&
0c&
0b&
1`&
0_&
1^&
0\&
0[&
1Y&
1X&
0W&
0U&
1T&
0S&
1R&
1Q&
0K&
1J&
0I&
0F&
1C&
1?&
0>&
1=&
1<&
0:&
09&
17&
15&
04&
13&
02&
0/&
0,&
0+&
0%&
0$&
1#&
1}%
1y%
0v%
1r%
0l%
0k%
1j%
0i%
0h%
0g%
1f%
0e%
1d%
1c%
1_%
0^%
0]%
1[%
0Z%
1Y%
0W%
0V%
1T%
1S%
0R%
0P%
1O%
0N%
1M%
1L%
1E%
1C%
1B%
1?%
1>%
1;%
1:%
18%
17%
13%
12%
10%
1.%
1,%
1+%
1(%
0"%
0!%
1}$
0|$
1z$
1y$
0x$
1s$
0p$
1n$
0i$
0h$
1f$
0e$
0b$
1a$
0`$
0^$
0]$
1\$
1X$
0U$
1T$
1L$
0K$
1J$
0I$
0G$
0F$
1E$
0C$
1=$
1<$
0:$
19$
07$
06$
15$
00$
1-$
0+$
1&$
1%$
0#$
1"$
0~#
0|#
0{#
0z#
0y#
0w#
0s#
0q#
0m#
0l#
0k#
0g#
0e#
0d#
0c#
0b#
0`#
0_#
0^#
0Z#
0Y#
1W#
0V#
1T#
1S#
0R#
1M#
0J#
1H#
0C#
0B#
1@#
0?#
07#
06#
15#
11#
1-#
0*#
1&#
0~"
0}"
1|"
0{"
0z"
1v"
1u"
0s"
1r"
0p"
0o"
1n"
0i"
1f"
0d"
1_"
1^"
0\"
1["
1X"
1V"
1S"
1R"
1O"
1N"
1K"
1H"
1G"
1F"
1C"
1A"
1?"
1<"
1;"
19"
18"
18(
1D(
1H(
1J(
0P(
1R(
1m8
1.*
1-*
0+*
1**
0(*
0'*
1&*
0!*
1|)
0z)
1u)
1t)
0r)
1q)
1U,
0P,
0O,
1M,
0L,
1J,
1I,
0H,
1C,
0@,
1>,
09,
08,
16,
05,
1'/
1&/
0$/
1#/
0!/
0~.
1}.
0x.
1u.
0s.
1n.
1m.
0k.
1j.
0Q/
1P/
0O/
0M/
0L/
1K/
1G/
0D/
1C/
1;/
0:/
19/
08/
06/
05/
14/
02/
0t/
0s/
1q/
0p/
1n/
1m/
0l/
1g/
0d/
1b/
0]/
0\/
1Z/
0Y/
1(2
1&2
1%2
1"2
1!2
1|1
1{1
1y1
1x1
1t1
1s1
1q1
1o1
1m1
1l1
1i1
1Q2
0O2
1N2
0M2
1L2
1K2
1G2
0F2
0E2
1C2
0B2
1A2
0?2
0>2
1<2
1;2
0:2
082
172
062
152
142
1O5
0M5
1L5
0K5
1J5
1I5
1E5
0D5
0C5
1A5
0@5
1?5
0=5
0<5
1:5
195
085
065
155
045
135
125
1m)
1k)
1h)
1g)
1d)
1c)
1`)
1])
1\)
1[)
1X)
1V)
1T)
1Q)
1P)
1N)
1M)
1L)
1K)
0J)
0(,
0',
1&,
1",
1|+
0y+
1u+
0o+
0n+
1m+
0l+
0k+
1j+
0y,
0w,
0v,
0u,
0t,
0r,
0n,
0l,
0h,
0g,
0f,
0b,
0`,
0_,
0^,
0],
0[,
0Z,
0Y,
1X,
0p2
0o2
1n2
1j2
1f2
0c2
1_2
0Y2
0X2
1W2
0V2
0U2
1T2
1)5
0'5
1&5
0%5
0"5
1}4
1y4
0x4
1w4
1v4
0t4
0s4
1q4
1o4
0n4
1m4
0l4
0i4
0f4
0e4
1d4
1#8
0"8
1!8
1|7
0y7
0u7
1t7
0s7
0r7
1p7
1o7
0m7
0k7
1j7
0i7
1h7
1e7
1b7
1a7
0`7
1r5
1p5
1m5
1l5
1i5
1h5
1e5
1b5
1a5
1`5
1]5
1[5
1Y5
1V5
1U5
1S5
0R5
0I8
0D8
0@8
1?8
1>8
0<8
1;8
188
178
068
058
048
138
128
0-8
0)8
0'8
1&8
157
127
007
1/7
0.7
1-7
0,7
1+7
1&7
1%7
0$7
1#7
1"7
1!7
1~6
1}6
1{6
1z6
0y6
1v6
0u6
1t6
0s6
0r6
1q6
1o6
1m6
0l6
0Y7
1X7
0W7
1V7
1T7
1Q7
0N7
1M7
1L7
0J7
0I7
0H7
1F7
1E7
0D7
1C7
0B7
1A7
0@7
1?7
1=7
0;7
1:7
154
144
134
004
1/4
0.4
0-4
1,4
0*4
0&4
0%4
1#4
0"4
1!4
1~3
0}3
1|3
1{3
0z3
1y3
0w3
1v3
0u3
1s3
1r3
1q3
1p3
0o3
1n3
0[4
1Z4
1X4
1V4
1U4
0T4
1R4
1O4
1N4
1M4
0K4
1J4
1G4
0F4
1C4
1A4
1?4
0=4
0<4
0:4
151
141
021
111
001
0/1
1*1
1)1
0'1
1&1
1!1
1~0
1}0
1{0
0y0
1x0
0w0
0v0
1s0
0]1
1Z1
0Y1
0X1
1W1
0T1
1S1
0P1
1O1
0N1
1K1
0I1
0H1
1C1
0B1
0A1
1@1
0=1
19.
05.
03.
0..
0-.
0,.
0(.
0|-
0z-
1x-
0w-
0v-
1u-
0t-
0s-
1r-
0\.
0[.
0X.
1V.
1U.
0L.
0E.
0D.
0B.
0A.
1@.
0?.
1A+
1?+
09+
07+
06+
05+
01+
00+
1(+
1~*
1}*
1|*
1`+
1_+
1\+
1[+
1X+
1U+
1T+
1P+
1I+
1H+
1E+
0B+
0$:
1{9
1z9
1y9
1x9
1w9
1t9
0p9
1n9
1k9
0j9
1d9
1b9
1a9
1`9
1I:
0C:
0B:
0?:
0<:
1::
19:
07:
06:
14:
03:
12:
0*:
0):
#91800
1"
1T!
b111010000111110001000100000000001101 N:
b100110000001000110010011001100000 O:
b1001001000011111000100010000000000111101 P:
b100100100000011000100110011001000000 Q:
b111000010010111111010111001100100110000 R:
b111001101000110001001100110011000100 S:
b1011111010110110110110001001100101011100 T:
b101010101001001110110011010100000 U:
b111010010110011011111011100110101011101 V:
b100101010101100000110011001010100000 W:
b11101000110100110100101111111011010100 X:
b10111001011000111010001000100010000 Y:
b10011110001110110001111101010110011101100 "F
b1010001100001001100000000101101000000000 #F
b1100111011111010011001100001101110100101000 $F
b100001000001000001100010011100010100000000000 %F
b11100101001101010111101111011011100001010100 &F
b1010010010101000010000101000010100000000 'F
b101010100110110001011000010110100101101011101000001000 xK
b1100100111101100001001010100010101000000 yK
b1111100100100011110100010001111011000110000000000000000 zK
b10000001000000001000100000000000000000000000000000 {K
b1110001101011100010101101001001111000100010001001000110010111100 HQ
b100010000011000010010110010000101001001010000100000000000000 IQ
b1111111010011000001010001110010110000000010110111011111000001 P!
b1111100111110010000000101001101001111011101011001000100011101100 Q!
b101011110011101100100100010110100111000010100010010001000 R!
b1111010001100010011010010101110000010110100101010000110010111100 S!
b10010110101010110101100000101101 H!
b101110010110000100100101011100 J!
b11110100000000000111101011101000 L!
b1111001001100000110100111110010 N!
b10110010101001110010011001100101 I!
b11011110100011100010100010111101 K!
b11100010110010100100111011000101 M!
b11100111011101101001011011001110 O!
1gY
1dY
1cY
0_Y
1^Y
0[Y
1ZY
0YY
1WY
1VY
0SY
1QY
1PY
0OY
1NY
1KY
0JY
1HY
1EY
0CY
1BY
0?Y
0=Y
0<Y
0;Y
07Y
06Y
14Y
12Y
1.Y
1-Y
1,Y
1+Y
1*Y
0b
1_
1^
1\
0Z
1Y
0W
0V
0U
0T
1S
0R
0P
1L
0K
0F
0E
1A
1;
0:
09
15
03
01
00
0/
1.
1-
0,
0*
0(
1&
0LN
0BN
1:N
09N
07N
16N
03N
01N
00N
0*N
0iM
0hM
0gM
1eM
0cM
1aM
0ZM
0YM
0UM
0TM
1QM
1PM
1OM
1NM
0MM
0HM
0FM
1CM
18M
16M
14M
02M
10M
0-M
1,M
1)M
0%M
1$M
1#M
0"M
1~L
1|L
0zL
0xL
1uL
0[L
0YL
0XL
0VL
1TL
0SL
1QL
0OL
0JL
1IL
0HL
0BL
0>L
0=L
1;L
19L
08L
15L
03L
12L
11L
1.L
0-L
1SJ
0RJ
1QJ
1LJ
0FJ
1EJ
0BJ
1@J
1>J
0=J
1<J
19J
08J
14J
1#J
1!J
1wI
0uI
1pI
1nI
0mI
1lI
1jI
1iI
0hI
0fI
1eI
0dI
1cI
1_I
0\I
0[I
1LI
1JI
0GI
1FI
1EI
1DI
1AI
1=I
1<I
16I
10I
1+I
0fG
0dG
0`G
0]G
1[G
1ZG
0YG
1XG
1WG
0TG
0SG
0PG
0OG
1MG
0KG
1EG
1DG
0CG
1AG
1@G
0?G
1<G
0;G
09G
01G
1-G
1+G
1*G
0)G
1(G
0%G
0~F
1}F
0{F
1yF
1tF
1sF
1mF
1\F
1YF
1WF
0VF
0UF
1SF
0RF
1QF
0NF
1MF
1KF
1EF
0CF
1BF
0?F
0>F
0=F
1:F
19F
07F
16F
05F
1"D
0zC
0yC
0vC
0sC
1qC
1pC
0nC
0mC
1kC
0jC
1iC
0aC
0`C
0VC
1OC
1NC
1MC
1LC
1KC
1HC
0DC
1BC
1?C
0>C
18C
16C
15C
14C
0.C
1-C
0,C
1+C
1)C
1&C
0#C
1"C
1!C
0}B
0|B
0{B
1yB
1xB
0wB
1vB
0uB
1tB
0sB
1rB
1pB
0nB
1mB
1eB
1bB
0`B
1_B
0^B
1]B
0\B
1[B
1VB
1UB
0TB
1SB
1RB
1QB
1PB
1OB
1MB
1LB
0KB
1HB
0GB
1FB
0EB
0DB
1CB
1AB
1?B
0>B
0.@
1-@
1+@
1)@
1(@
0'@
1%@
1"@
1!@
1~?
0|?
1{?
1x?
0w?
1t?
1r?
1p?
0n?
0m?
0k?
1`?
1_?
1^?
0[?
1Z?
0Y?
0X?
1W?
0U?
0Q?
0P?
1N?
0M?
1L?
1K?
0J?
1I?
1H?
0G?
1F?
0D?
1C?
0B?
1@?
1??
1>?
1=?
0<?
1;?
04?
11?
00?
0/?
1.?
0+?
1*?
0'?
1&?
0%?
1"?
0~>
0}>
1x>
0w>
0v>
1u>
0r>
1d>
1c>
0a>
1`>
0_>
0^>
1Y>
1X>
0V>
1U>
1P>
1O>
1N>
1L>
0J>
1I>
0H>
0G>
1D>
0?<
0><
0;<
19<
18<
0/<
0(<
0'<
0%<
0$<
1#<
0"<
1x;
0t;
0r;
0m;
0l;
0k;
0g;
0];
0[;
1Y;
0X;
0W;
1V;
0U;
0T;
1S;
1K;
1J;
1G;
1F;
1C;
1@;
1?;
1;;
14;
13;
10;
0-;
1&;
1$;
0|:
0z:
0y:
0x:
0t:
0s:
1k:
1c:
1b:
1a:
1NR
1LR
1HR
1GR
0FR
0BR
0@R
0>R
0<R
08R
15R
11R
10R
1,R
1+R
0*R
1A=
1?=
09=
07=
01=
00=
1(=
0"=
1~<
1}<
1|<
0{<
1uR
0qR
0nR
0kR
0jR
0dR
1_R
0ZR
0WR
0VR
0QR
1PR
0.>
0+>
1)>
1(>
0v=
0r=
1q=
0p=
1rS
1oS
0kS
0hS
0fS
0bS
0_S
0^S
0ZS
1XS
1TS
0RS
1QS
15A
02A
11A
00A
0/A
1+A
1*A
0)A
1(A
0'A
1&A
0"A
0!A
1}@
1{@
0y@
1x@
0w@
0v@
0s@
0q@
1?T
1>T
1=T
0<T
0;T
0:T
08T
15T
04T
13T
0.T
1-T
1*T
0)T
1&T
1%T
0$T
0#T
0!T
0~S
1}S
1zS
1xS
0.B
1)B
0'B
1"B
1!B
1~A
0|A
1xA
1tA
1rA
0kA
1EU
1BU
0<U
18U
16U
12U
1*U
1)U
0%U
1#U
0"U
1}T
0|T
1'E
1$E
0"E
1!E
0~D
1}D
0|D
1{D
1vD
1uD
1tD
1sD
1rD
1qD
1mD
1lD
0kD
1hD
0gD
1fD
1eD
0dD
1cD
1aD
1_D
1^D
0hU
1fU
1aU
0^U
1]U
1\U
0ZU
0YU
0WU
0SU
0OU
0JU
0HU
0nE
1EH
1BH
1AH
1@H
0>H
0<H
08H
17H
05H
03H
12H
11H
1/H
0.H
1)H
1'H
0&H
0%H
1$H
0#H
1"H
1~G
1{G
0zG
1xG
1wG
0vG
1sG
0rG
0pG
0xH
0vH
1sH
1qH
0pH
1oH
0nH
1kH
1jH
0iH
1eH
0dH
0cH
1bH
0`H
0_H
0^H
1]H
1\H
0[H
1ZH
0WH
1VH
15K
11K
00K
0/K
1.K
1-K
1,K
0+K
1)K
0'K
0&K
1"K
1~J
1}J
1zJ
0xJ
0vJ
0rJ
1pJ
0lJ
1jK
1fK
1aK
1]K
1\K
0VK
1UK
1PK
1NK
0MK
1LK
1KK
0"W
0~V
0}V
0xV
0wV
1vV
1uV
0tV
0sV
1pV
1nV
0mV
1lV
1hV
0fV
0eV
1bV
0aV
1`V
0_V
0^V
0XV
1WV
1VV
1SV
0RV
1>Q
1;Q
13Q
00Q
0+Q
1)Q
0'Q
1%Q
0"Q
1}P
0{P
1zP
1yP
1vP
1uP
1tP
0OW
0NW
0MW
0LW
1JW
0HW
1FW
1EW
0?W
0>W
1=W
1<W
15W
02W
0+W
1(W
0nO
0[O
0SO
0RO
0LO
1[P
1XP
1PP
0MP
0HP
1FP
0DP
1BP
0?P
1<P
0:P
19P
18P
15P
14P
13P
0DX
0BX
0AX
0<X
0;X
1:X
19X
08X
07X
14X
12X
1/X
0.X
0)X
0(X
0'X
1&X
1%X
0$X
1#X
1"X
0!X
0~W
0}W
1|W
0zW
0yW
0xW
1tW
0rW
0kW
1hW
1<Q
0;Q
0:Q
18Q
05Q
03Q
1+Q
0$Q
0zP
0uP
1XD
1UD
0SD
1RD
0QD
1PD
0OD
1ND
1ID
1HD
1GD
1FD
1ED
1DD
1@D
1?D
0>D
1;D
0:D
19D
18D
07D
16D
14D
12D
11D
1?V
1<V
04V
02V
10V
0/V
0+V
0*V
0(V
0'V
0%V
0$V
0#V
0!V
0}U
1zU
0wU
0tU
0'E
0$E
1xD
0eD
0bD
0_D
0^D
1c@
0`@
1_@
0^@
0]@
1Y@
1X@
0W@
1V@
0U@
1T@
0P@
0O@
1M@
1K@
0I@
1H@
0G@
0F@
0C@
0A@
1rT
1oT
1nT
1mT
1lT
0jT
0iT
0hT
0gT
1fT
1dT
0cT
1_T
1^T
1]T
0\T
0ZT
1YT
1UT
1ST
1QT
1PT
0OT
1NT
1KT
1IT
05A
1.A
0+A
1)A
1"A
1!A
1u@
1s@
1s<
1q<
0k<
0i<
0c<
0b<
1Z<
0T<
1R<
1Q<
1P<
0O<
1FS
0DS
1BS
0@S
0?S
1;S
1:S
07S
16S
14S
01S
10S
0-S
0,S
0)S
0(S
1'S
0"S
0|R
1{R
0A=
1;=
1:=
13=
0(=
1$=
1#=
0}<
0s<
1m<
1l<
1e<
0Z<
1V<
1U<
0Q<
1l=
1k=
0j=
0i=
1h=
0f=
0e=
1c=
1`=
0]=
1\=
0[=
0W=
1V=
0S=
0O=
0N=
1M=
1L=
0J=
0I=
0G=
0D=
1C=
16>
00>
0->
0)>
1~=
0w=
1u=
1t=
0c@
1\@
0Y@
1W@
1P@
1O@
1E@
1C@
1dA
0cA
1aA
0]A
0\A
1[A
0ZA
1WA
0TA
1QA
1NA
1MA
0LA
0IA
0HA
0FA
1EA
0BA
1@A
1=A
1;A
14B
10B
1-B
0,B
1+B
0(B
1'B
0&B
1%B
0"B
0!B
0~A
0}A
1{A
1zA
1wA
0vA
0tA
0rA
1qA
0XD
0UD
1KD
08D
05D
02D
01D
1SE
1RE
1PE
0OE
0ME
1LE
1KE
1JE
1IE
0FE
0DE
1BE
0AE
0@E
0<E
0;E
0:E
07E
14E
02E
11E
1.E
0-E
1,E
1+E
0*E
1{E
0wE
0uE
1tE
1mE
1lE
1hE
1fE
1eE
0`E
1_E
1^E
0]E
1\E
1YE
1VE
1YP
0XP
0WP
1UP
0RP
0PP
1HP
0AP
09P
04P
0AO
0?O
0>O
08O
17O
15O
04O
01O
1/O
1.O
1,O
0%O
0#O
1!O
0}N
1|N
0zN
1yN
0xN
0wN
1tN
1pN
0hN
1eN
1vO
0uO
1qO
0kO
0fO
1cO
0aO
1`O
1_O
0^O
0]O
1\O
1ZO
1SO
07O
16O
05O
13O
10O
0.O
1&O
1}N
0uN
0pN
1wO
0vO
0pO
0_O
0RE
1OE
1EE
12E
0/E
0,E
0+E
0{E
0^E
1cA
1\A
0YA
0WA
0PA
0OA
0EA
0CA
04B
1(B
1!B
1~A
1tA
1rA
0k=
1e=
1d=
1]=
0R=
1N=
0M=
1I=
1x=
0t=
#93600
b10110001111011110110001001100011 d
b101011100111000011100001010 e
0"
0)Y
1(Y
0'Y
1&Y
0$Y
0#Y
1!Y
0zX
1xX
0uX
1sX
1qX
0pX
1oX
0nX
1mX
0kX
0jX
0hX
0u!
1t!
0s!
1r!
0p!
0o!
1m!
0h!
1f!
0c!
1a!
1_!
0^!
1]!
0\!
1[!
0Y!
0X!
0V!
1fX
0eX
0dX
1aX
1^X
0\X
0[X
1ZX
1UX
1QX
1OX
0NX
0MX
1JX
0G!
1F!
1E!
1D!
1C!
0?!
0>!
1<!
0;!
0:!
09!
06!
15!
04!
13!
12!
10!
1/!
0*!
1)!
0(!
1'!
1&!
0$!
0#!
1!!
0}
1|
0{
1y
1x
1w
0u
1s
0n
0m
1h
1g
1f
0T!
0r(
1q(
0p(
1o(
0m(
0l(
1j(
0e(
1c(
0`(
1^(
1\(
0[(
1Z(
0Y(
1X(
0V(
0U(
0S(
16"
05"
04"
11"
1."
0,"
0+"
1*"
1%"
1!"
1}!
0|!
0{!
1x!
b1 vQ
b0 pQ
b0 mQ
b0 gQ
b1 ^Q
b1 XQ
b0 [Q
b1 LQ
b0 OQ
0SQ
1VQ
0YQ
1bQ
0eQ
0kQ
1tQ
0zQ
b111111010100011000111100011110101 KQ
b101011100111000011100001010 NQ
b111110101000110001111000111101011 QQ
b1010111001110000111000010100 TQ
b111110101000110001111000111101011 WQ
b101011100111000011100001010 ZQ
b111110101000110001111000111101011 ]Q
b1010111001110000111000010100 `Q
b111111010100011000111100011110101 cQ
b0 fQ
b111111010100011000111100011110101 iQ
b0 lQ
b1010111001110000111000010100 oQ
b0 rQ
b111111010100011000111100011110101 uQ
b111111010100011000111100011110101 xQ
0#)
1")
0!)
1|(
0{(
0y(
1v(
0t(
1k'
1j'
0i'
0h'
1f'
1c'
0b'
0a'
1_'
1^'
0]'
0\'
1T'
1S'
1Q'
1L'
1I'
0G'
0F'
1E'
1D'
1B'
0@'
0?'
1='
0;'
15'
12'
0.'
0,'
0)'
0('
0%'
0$'
0!'
0|&
0{&
0z&
0w&
0u&
0s&
0p&
0o&
0m&
0k&
1j&
0i&
0e&
0d&
1c&
1b&
0`&
0^&
0]&
1\&
1[&
1Z&
0Y&
0X&
1W&
1U&
0T&
1S&
0R&
0N&
0J&
0H&
0G&
0D&
0C&
0@&
0?&
0=&
0<&
08&
07&
05&
03&
01&
00&
0-&
1*&
0)&
1(&
0'&
1%&
1$&
0"&
1{%
0y%
1v%
0t%
0r%
1q%
0p%
1o%
0n%
1l%
1k%
1i%
1h%
0f%
0d%
0c%
0`%
0_%
0\%
0[%
0Y%
0X%
0T%
0S%
0Q%
0O%
0M%
0L%
0I%
1F%
0E%
1D%
0C%
1A%
1@%
0>%
19%
07%
14%
02%
00%
1/%
0.%
1-%
0,%
1*%
1)%
1'%
1&%
0%%
1!%
0~$
0}$
1x$
0v$
1m$
1h$
0g$
0f$
0d$
0c$
1b$
1]$
1Z$
0X$
0W$
1V$
1U$
1S$
0Q$
0P$
1N$
0L$
1F$
1C$
0A$
1@$
0?$
1>$
0=$
0<$
17$
05$
04$
10$
1+$
0*$
1)$
0($
1'$
0&$
0%$
0"$
1~#
1}#
1{#
1y#
1x#
1w#
1v#
1r#
1q#
1p#
1o#
1k#
1j#
1f#
1d#
1b#
1a#
1`#
1_#
1^#
0]#
1Y#
0X#
0W#
1R#
0P#
1G#
1B#
0A#
0@#
0>#
0=#
1<#
08#
17#
16#
01#
1/#
0&#
0!#
1~"
1}"
1{"
1z"
0u"
0r"
1p"
1o"
0n"
0m"
0k"
1i"
1h"
0f"
1d"
0^"
0["
1T"
1Q"
0O"
0N"
1M"
1L"
1J"
0H"
0G"
1E"
0C"
1="
1:"
06(
14(
0>(
1<(
1@(
0F(
0J(
0L(
1P(
1i)
1f)
0d)
0c)
1b)
1a)
1_)
0])
0\)
1Z)
0X)
1R)
1O)
13*
0-*
0**
1(*
1'*
0&*
0%*
0#*
1!*
1~)
0|)
1z)
0t)
0q)
1-/
0+/
1*/
0)/
1(/
0'/
0&/
1!/
0}.
0|.
1x.
1s.
0r.
1q.
0p.
1o.
0n.
0m.
0j.
0S/
1Q/
1L/
1I/
0G/
0F/
1E/
1D/
1B/
0@/
0?/
1=/
0;/
15/
12/
0N2
0L2
0K2
0H2
0G2
0D2
0C2
0A2
0@2
0<2
0;2
092
072
052
042
012
0&5
0$5
0#5
0~4
0}4
0z4
0y4
0w4
0v4
0r4
0q4
0o4
0m4
0k4
0j4
0g4
0O5
0L5
1K5
0J5
0F5
0E5
1D5
1C5
0A5
0?5
0>5
1=5
1<5
1;5
0:5
095
185
165
055
145
035
0/5
1}7
1z7
0x7
0w7
1v7
1u7
1s7
0q7
0p7
1n7
0l7
1f7
1c7
1I8
1A8
1@8
0?8
0>8
1<8
198
088
078
158
148
038
028
1*8
1)8
1'8
0&8
0u5
0r5
0p5
0m5
0l5
0i5
0h5
0e5
0b5
0a5
0`5
0]5
0[5
0Y5
0V5
0U5
0S5
1R5
0w2
1u2
0t2
1s2
0r2
1p2
1o2
0m2
1h2
0f2
1c2
0a2
0_2
1^2
0]2
1\2
0[2
1Y2
1X2
1V2
1U2
0T2
1)2
0(2
1'2
0&2
1$2
1#2
0!2
1z1
0x1
1u1
0s1
0q1
1p1
0o1
1n1
0m1
1k1
1j1
1h1
1g1
0f1
1y/
0w/
1s/
0r/
0q/
1l/
0j/
1a/
1\/
0[/
0Z/
0X/
0W/
1V/
1y,
1x,
1v,
1t,
1s,
1r,
1q,
1m,
1l,
1k,
1j,
1f,
1e,
1a,
1_,
1],
1\,
1[,
1Z,
1Y,
0X,
0S,
1O,
0N,
0M,
1H,
0F,
1=,
18,
07,
06,
04,
03,
12,
0/,
1-,
0),
1(,
1',
0",
1~+
0u+
0p+
1o+
1n+
1l+
1k+
0j+
0;.
09.
07.
11.
10.
1/.
1-.
1*.
1).
1(.
0'.
1&.
0#.
0".
1|-
1v-
1s-
0r-
1a.
1\.
1[.
0Y.
1T.
0R.
1O.
1J.
1I.
0F.
1E.
1D.
1A.
0@.
1>.
0%:
0!:
0|9
0{9
0w9
0v9
1u9
0q9
1p9
0o9
1m9
1l9
0h9
1e9
0d9
1c9
0a9
0`9
1K:
1G:
1D:
1C:
0A:
1?:
1>:
0::
17:
05:
04:
10:
1,:
1):
037
027
017
0+7
0*7
1(7
0%7
0#7
0"7
0{6
1y6
1x6
0w6
0q6
1p6
0o6
0m6
1l6
0X7
0V7
0T7
0Q7
0P7
0M7
0L7
0F7
0E7
0C7
0A7
0?7
0=7
0:7
054
044
014
104
0/4
1.4
1-4
1)4
1'4
1&4
1%4
0#4
1"4
0!4
0~3
1}3
0|3
0{3
1z3
0y3
0x3
1w3
0v3
1u3
0t3
0s3
0p3
1o3
0n3
1]4
0Z4
1Y4
0X4
1W4
0V4
0U4
0Q4
0O4
0N4
0M4
1K4
0J4
0G4
1F4
0E4
0C4
1B4
0A4
1@4
0?4
1>4
1=4
1:4
191
161
051
041
121
101
1/1
0.1
0-1
0)1
0&1
0$1
0#1
0~0
1|0
1z0
1y0
1w0
1u0
0r0
0q0
1p0
0_1
1]1
1\1
0[1
0Z1
1U1
0S1
0R1
1Q1
1P1
1N1
1I1
0F1
1E1
0D1
0C1
0?1
0A+
1=+
1;+
1:+
17+
14+
10+
0/+
0*+
1&+
1$+
1#+
1!+
1e+
0_+
0\+
0[+
1Z+
1Y+
0X+
0U+
0T+
1S+
1R+
0P+
1N+
0H+
0E+
#95400
1"
1T!
b111111101111010000100110010011011100 N:
b10000100011000001100000100001 O:
b101101000111100001011110101110000101000 P:
b10010111000110011100001110001111000100 Q:
b1001010111111101100000101000011110001001 R:
b101000010001110011110001110000110000 S:
b101100101001001001011111101111010010000 T:
b10011010100010000100000010000101000100 U:
b1010100010101110011100001110000101000001 V:
b0 W:
b110100010111101000110011100010010000 X:
b1011111101000010101011100011101010100 Y:
b100001100101010000010111011011111110110001 "F
b100010010001011100000100000000000001000 #F
b1011110001001001001100101000000011010110111000 $F
b1110100110110011010101110101001000000000 %F
b11000010011111000100001100110101111110011101 &F
b101110100100101110110011001000100000000000 'F
b110011101111010100101010101111000110011000011101100 xK
b10101011000110010000111001010110000000000 yK
b1111000110000001011101111001001110111001000100000000000 zK
b10000110101000010000101100010000100010000000000000 {K
b1111000101011100011000010011011010100100110110010010010010001000 HQ
b100000000001000010101000100100001000000001000001000000000000 IQ
b1111111001010110011100100100011101010001101101010000110011011110 P!
b1111111010011000001010001110010110000000010110111011111000001 Q!
b1111100111110010000000101001101001111011101011001000100011101100 R!
b101011110011101100100100010110100111000010100010010001000 S!
b10110001111011110110001001100011 H!
b10010110101010110101100000101101 J!
b101110010110000100100101011100 L!
b11110100000000000111101011101000 N!
b101011100111000011100001010 I!
b10110010101001110010011001100101 K!
b11011110100011100010100010111101 M!
b11100010110010100100111011000101 O!
1iY
0gY
0fY
0dY
1aY
1`Y
1_Y
0^Y
1]Y
1\Y
1[Y
0ZY
1YY
1XY
0WY
0TY
0RY
0QY
0PY
0NY
0KY
1JY
0HY
1GY
0BY
1AY
0@Y
1?Y
19Y
04Y
10Y
1/Y
0,Y
0+Y
0*Y
0a
0_
0^
0X
1U
0Q
0O
1N
1M
0J
1F
1D
0A
0?
0;
1:
19
08
17
11
10
1/
0.
1+
0)
0'
0&
0%
0$
1JN
1FN
1AN
1=N
1<N
06N
15N
10N
1.N
0-N
1,N
1+N
1kM
1gM
0fM
0eM
1dM
1cM
1bM
0aM
1_M
0]M
0\M
1XM
1VM
1UM
1RM
0PM
0NM
0JM
1HM
0DM
08M
06M
13M
11M
00M
1/M
0.M
1+M
1*M
0)M
1%M
0$M
0#M
1"M
0~L
0}L
0|L
1{L
1zL
0yL
1xL
0uL
1tL
1[L
1XL
1WL
1VL
0TL
0RL
0NL
1ML
0KL
0IL
1HL
1GL
1EL
0DL
1?L
1=L
0<L
0;L
1:L
09L
18L
16L
13L
02L
10L
1/L
0.L
1+L
0*L
0(L
0SJ
0QJ
1PJ
0JJ
1IJ
1HJ
1DJ
1BJ
1AJ
0<J
1;J
09J
18J
15J
12J
1%J
1"J
0}I
1|I
1{I
1zI
1yI
0vI
1uI
0tI
1rI
0qI
0pI
0lI
0kI
0jI
0gI
1dI
1aI
0_I
1^I
0]I
0ZI
1NI
0LI
1KI
0JI
1II
1GI
0DI
1CI
1?I
1>I
0=I
0<I
1;I
1:I
18I
17I
06I
14I
12I
11I
0+I
1bG
1_G
0[G
1YG
0XG
0WG
0RG
1OG
0NG
0MG
1LG
1KG
0JG
0GG
0FG
0DG
0AG
0@G
1>G
1;G
19G
13G
0-G
0+G
0*G
0(G
1%G
1{F
1uF
0tF
0sF
1rF
0oF
1nF
0mF
1^F
0\F
0[F
1ZF
0XF
1VF
1UF
1RF
1NF
0MF
0IF
1HF
0EF
0DF
0AF
1>F
0<F
09F
06F
15F
1$D
1~C
1{C
1zC
0xC
1vC
1uC
0qC
1nC
0lC
0kC
1gC
1cC
1`C
0WC
0SC
0PC
0OC
0KC
0JC
1IC
0EC
1DC
0CC
1AC
1@C
0<C
19C
08C
17C
05C
04C
0-C
0+C
0)C
0&C
0%C
0"C
0!C
0yB
0xB
0vB
0tB
0rB
0pB
0mB
0cB
0bB
0aB
0[B
0ZB
1XB
0UB
0SB
0RB
0MB
1KB
1JB
0IB
0CB
1BB
0AB
0?B
1>B
10@
0-@
1,@
0+@
1*@
0)@
0(@
0$@
0"@
0!@
0~?
1|?
0{?
0x?
1w?
0v?
0t?
1s?
0r?
1q?
0p?
1o?
1n?
1k?
0`?
0_?
0\?
1[?
0Z?
1Y?
1X?
1T?
1R?
1Q?
1P?
0N?
1M?
0L?
0K?
1J?
0I?
0H?
1G?
0F?
0E?
1D?
0C?
1B?
0A?
0@?
0=?
1<?
0;?
06?
14?
13?
02?
01?
1,?
0*?
0)?
1(?
1'?
1%?
1~>
0{>
1z>
0y>
0x>
0t>
1h>
1e>
0d>
0c>
1a>
1_>
1^>
0]>
0\>
0X>
0U>
0S>
0R>
0O>
1M>
1K>
1J>
1H>
1F>
0C>
0B>
1A>
1D<
1?<
1><
0<<
17<
05<
12<
1-<
1,<
0)<
1(<
1'<
1$<
0#<
1!<
0z;
0x;
0v;
1p;
1o;
1n;
1l;
1i;
1h;
1g;
0f;
1e;
0b;
0a;
1];
1W;
1T;
0S;
1P;
0J;
0G;
0F;
1E;
1D;
0C;
0@;
0?;
1>;
1=;
0;;
19;
03;
00;
0&;
1";
1~:
1}:
1z:
1w:
1s:
0r:
0m:
1i:
1g:
1f:
1d:
0NR
1MR
1JR
0HR
0CR
1BR
1@R
1;R
1:R
18R
07R
06R
13R
01R
1.R
1-R
0?=
1==
0;=
14=
0/=
1*=
0'=
1&=
1"=
1!=
0wR
0uR
0tR
0sR
1oR
1nR
0mR
1kR
0iR
0gR
1fR
1dR
0cR
0_R
0^R
0]R
0\R
1ZR
0YR
1XR
1WR
1SR
0PR
1z=
1v=
1r=
0q=
1o=
1vS
0rS
1pS
1nS
1mS
1lS
1kS
1jS
1iS
1gS
0eS
1dS
1cS
1bS
0aS
0`S
1[S
1ZS
1WS
1VS
0TS
0SS
0QS
0PS
1OS
19A
10A
1/A
0.A
0-A
0)A
0&A
1#A
0}@
1|@
1z@
1y@
1w@
0u@
0t@
0r@
1q@
1p@
0?T
16T
03T
12T
11T
1.T
0-T
0*T
1)T
0%T
0|S
0zS
0xS
0-B
1,B
0+B
1*B
1|A
0{A
0xA
1sA
0pA
1kA
0CU
0BU
0AU
1?U
1=U
0:U
17U
05U
04U
02U
1,U
1+U
0)U
1(U
1&U
0$U
0#U
1"U
0}T
1|T
0{D
0vD
0uD
0sD
0qD
0pD
1oD
0mD
1kD
1jD
0iD
1bD
0aD
1_D
1^D
0iU
1hU
0eU
0dU
1bU
0`U
1^U
0]U
0VU
0UU
0TU
1SU
1QU
0NU
1MU
0KU
1JU
0GU
1vE
1rE
1oE
1nE
1jE
0eE
0_E
1[E
1WE
1GH
0EH
0DH
0AH
1?H
1>H
1=H
0;H
0:H
07H
06H
15H
14H
00H
1.H
0+H
1*H
1(H
0'H
1%H
1#H
0"H
1!H
0}G
0|G
0{G
0xG
0wG
1uG
1rG
1pG
1zH
0tH
1rH
1nH
0kH
0eH
0aH
1^H
0]H
0\H
1[H
0ZH
0XH
0VH
1UH
17K
14K
13K
10K
1/K
0.K
0,K
1+K
0*K
0)K
0%K
1#K
0~J
0}J
1|J
0{J
0zJ
0wJ
1tJ
1sJ
1qJ
0pJ
1nJ
1mJ
1lJ
0jJ
0iJ
0jK
1iK
0fK
1eK
1cK
1`K
1^K
0]K
1[K
0ZK
1XK
1WK
0UK
1TK
1RK
1QK
0LK
0FK
1BK
1"W
1}V
1|V
1wV
0vV
1tV
1qV
0pV
1jV
0iV
0hV
0gV
1fV
1eV
0dV
0cV
0[V
1ZV
0YV
1XV
0WV
1UV
1TV
0SV
1PV
0OV
0MV
1EQ
1BQ
1AQ
0>Q
0<Q
08Q
17Q
13Q
12Q
1/Q
0.Q
0-Q
1,Q
0)Q
1'Q
0&Q
0%Q
1$Q
0#Q
1"Q
1~P
1|P
1{P
1xP
1wP
0vP
0tP
1sP
0pP
1PW
1MW
1LW
0KW
0JW
1HW
1GW
0FW
0BW
0AW
0@W
1?W
0=W
1;W
1:W
09W
08W
17W
05W
11W
00W
1.W
1-W
1)W
1^O
0XO
1WO
1RO
1NO
1MO
1bP
1_P
1^P
0[P
0YP
0UP
1TP
1PP
1OP
1LP
0KP
0JP
1IP
0FP
1DP
0CP
0BP
1AP
0@P
1?P
1=P
1;P
1:P
17P
16P
05P
03P
12P
0/P
1DX
1AX
1@X
1;X
0:X
18X
15X
04X
02X
0/X
0+X
1'X
1$X
0#X
0"X
1!X
0|W
1xW
0vW
1rW
0pW
1oW
1nW
1mW
1iW
0EQ
0BQ
0AQ
1;Q
06Q
1-Q
0,Q
1*Q
1)Q
0(Q
0sP
0ND
0ID
0HD
0FD
0DD
0CD
1BD
0@D
1>D
1=D
0<D
15D
04D
12D
11D
0=V
0<V
0;V
19V
16V
14V
03V
12V
11V
00V
1/V
1+V
0&V
1%V
1$V
1!V
0~U
1}U
0|U
0{U
1yU
0sU
0!E
0}D
0wD
0tD
0rD
0lD
0kD
0cD
0bD
0_D
0^D
1g@
1^@
1]@
0\@
0[@
0W@
0T@
1Q@
0M@
1L@
1J@
1I@
1G@
0E@
0D@
0B@
1A@
1@@
1vT
0rT
1pT
0mT
0lT
1kT
1jT
1iT
1gT
0dT
1cT
0]T
1\T
1[T
1ZT
0YT
0XT
1WT
0VT
0ST
0QT
0PT
1OT
0MT
0KT
0IT
09A
01A
00A
1,A
1'A
1%A
0$A
0#A
0{@
0x@
0w@
1u@
0q@
0p@
0q<
1o<
0m<
1f<
0a<
1\<
0Y<
1X<
1T<
1S<
0FS
1ES
1DS
0AS
0<S
06S
04S
02S
11S
0/S
1.S
1,S
0*S
0'S
0$S
1~R
0{R
0==
1;=
15=
1.=
1-=
0+=
0*=
1)=
0&=
0!=
0~<
0o<
1m<
1g<
1`<
1_<
0]<
0\<
1[<
0X<
0S<
0R<
0l=
1k=
1j=
1i=
0e=
0b=
1^=
0\=
0Z=
0Y=
0X=
1W=
1U=
1R=
1Q=
1M=
0L=
1K=
1J=
1F=
0C=
06>
14>
1/>
1)>
1'>
0|=
1{=
0x=
1w=
0g@
0_@
0^@
1Z@
1U@
1S@
0R@
0Q@
0K@
0H@
0G@
1E@
0A@
0@@
1hA
1gA
0dA
1bA
1_A
1YA
1WA
1VA
1UA
1TA
0QA
1OA
0NA
1KA
1HA
0GA
0DA
1CA
0@A
0?A
0=A
0;A
1.B
0,B
0*B
0(B
0'B
0%B
1"B
0~A
1}A
0|A
1{A
0zA
1xA
1vA
0tA
0rA
1pA
1oA
1nA
0RD
0PD
0JD
0GD
0ED
0?D
0>D
06D
05D
02D
01D
0QE
0PE
0OE
1ME
0JE
0GE
1FE
0EE
1DE
0BE
1@E
0?E
0>E
1=E
1<E
09E
17E
16E
05E
04E
03E
02E
01E
0.E
1,E
1+E
0)E
0tE
0rE
1qE
0oE
0lE
1kE
0iE
1eE
0bE
1aE
1_E
1]E
0bP
0_P
0^P
1XP
0SP
1JP
0IP
1GP
1FP
0EP
02P
1AO
0@O
1>O
0<O
09O
18O
15O
03O
11O
0/O
1.O
0-O
0,O
1*O
0)O
1'O
0"O
1{N
1wN
1vN
1uN
1rN
1qN
0nN
0mN
1lN
1jN
1fN
1"P
1}O
1|O
0wO
1rO
0qO
1mO
1lO
1bO
0`O
1_O
0^O
0WO
0SO
1PO
0NO
0MO
0HO
1@O
1=O
1<O
06O
01O
1(O
0'O
1%O
0$O
1#O
1nN
0"P
0}O
0|O
1vO
1dO
0cO
0PO
0LE
1JE
0DE
1AE
1?E
19E
18E
10E
1/E
0,E
0+E
0vE
0mE
0kE
0eE
0dE
0\E
0[E
0gA
0_A
0^A
1ZA
0UA
0SA
1RA
1QA
0KA
0HA
1GA
1EA
1AA
1@A
1&B
1$B
0#B
0"B
0vA
0pA
0oA
0g=
1e=
0_=
1X=
0W=
0U=
1T=
1S=
0P=
0K=
0J=
1,>
1$>
0!>
#97200
b11000000001110110010001010000000 d
b10000011001000010000100100000 e
0"
0(Y
0&Y
1$Y
0~X
0}X
1zX
0xX
0wX
0vX
1uX
0sX
0oX
0mX
1kX
0t!
0r!
1p!
0l!
0k!
1h!
0f!
0e!
0d!
1c!
0a!
0]!
0[!
1Y!
0gX
0fX
0bX
0aX
1`X
0YX
0UX
1SX
0QX
0PX
0OX
0KX
0JX
1IX
0F!
0E!
0D!
0C!
0A!
0@!
0=!
0<!
1;!
19!
18!
07!
16!
02!
11!
0/!
0+!
1*!
0)!
0&!
0%!
0!!
1}
0|
0y
0x
1v
0s
1r
0q
1p
1n
1m
0k
0T!
0q(
0o(
1m(
0i(
0h(
1e(
0c(
0b(
0a(
1`(
0^(
0Z(
0X(
1V(
07"
06"
02"
01"
10"
0)"
0%"
1#"
0!"
0~!
0}!
0y!
0x!
1w!
1wQ
b0 vQ
1kQ
b0 jQ
0hQ
b1 gQ
1SQ
b0 RQ
0VQ
b1 UQ
1MQ
b0 LQ
b0 KQ
b0 NQ
b0 QQ
b111011111001101111011110110111111 TQ
b111101111100110111101111011011111 WQ
b10000011001000010000100100000 ZQ
b111011111001101111011110110111111 ]Q
b10000011001000010000100100000 `Q
b111101111100110111101111011011111 cQ
b111101111100110111101111011011111 fQ
b0 iQ
b10000011001000010000100100000 lQ
b0 oQ
b0 uQ
b111101111100110111101111011011111 xQ
1u(
1y(
0z(
1#)
0")
1%)
1p'
1n'
0l'
1h'
1g'
0d'
1b'
1a'
1`'
0_'
1]'
1Y'
1W'
0U'
0P'
0N'
0L'
0K'
0J'
0I'
0E'
0D'
0C'
0B'
0>'
0='
09'
07'
05'
04'
03'
02'
01'
00'
0j&
0h&
0c&
0b&
0a&
0\&
0[&
0Z&
0W&
0V&
0U&
0S&
0Q&
1F&
1C&
1>&
19&
16&
15&
1/&
0*&
0(&
0&&
0%&
0$&
0#&
0}%
0|%
0{%
0z%
0v%
0u%
0q%
0o%
0m%
0l%
0k%
0j%
0i%
0h%
1g%
1f%
1e%
1d%
1c%
1a%
1`%
1^%
1]%
1\%
1[%
1Y%
1X%
1W%
1V%
1T%
1S%
1P%
1O%
1N%
1M%
1L%
1J%
1I%
1H%
1G%
1E%
1C%
0A%
1=%
1<%
09%
17%
16%
15%
04%
12%
1.%
1,%
0*%
0#%
0!%
1~$
1{$
0z$
0y$
0x$
1v$
0s$
0r$
0l$
0j$
0h$
1g$
1`$
1^$
0\$
1X$
1W$
0T$
1R$
1Q$
1P$
0O$
1M$
1I$
1G$
0E$
0@$
0>$
1<$
08$
07$
14$
02$
01$
00$
1/$
0-$
0)$
0'$
1%$
1|#
1z#
0y#
0v#
1u#
1t#
1s#
0q#
1n#
1m#
1g#
1e#
1c#
0b#
1]#
1\#
1Z#
1X#
1V#
1U#
0T#
1Q#
1P#
1N#
1I#
0G#
0F#
1E#
1C#
1A#
1?#
1>#
1=#
0<#
0;#
09#
07#
06#
05#
04#
00#
0/#
0.#
0-#
0)#
0(#
0$#
0"#
0~"
0}"
0|"
0{"
0z"
0x"
0v"
0q"
0p"
0o"
0j"
0i"
0h"
0e"
0d"
0c"
0a"
0_"
0X"
0V"
0T"
0S"
0R"
0Q"
0M"
0L"
0K"
0J"
0F"
0E"
0A"
0?"
0="
0<"
0;"
0:"
09"
08"
04(
1:(
08(
1F(
0H(
0P(
03*
00*
0.*
0)*
0(*
0'*
0"*
0!*
0~)
0{)
0z)
0y)
0w)
0u)
1{,
1w,
1u,
0t,
0q,
1p,
1o,
1n,
0l,
1i,
1h,
1b,
1`,
1^,
0],
0*/
0(/
1&/
0"/
0!/
1|.
0z.
0y.
0x.
1w.
0u.
0q.
0o.
1m.
1O/
1M/
0K/
1G/
1F/
0C/
1A/
1@/
1?/
0>/
1</
18/
16/
04/
0u/
0s/
1r/
1o/
0n/
0m/
0l/
1j/
0g/
0f/
0`/
0^/
0\/
1[/
1(2
1&2
0$2
1~1
1}1
0z1
1x1
1w1
1v1
0u1
1s1
1o1
1m1
0k1
0)5
1"5
1}4
1x4
1s4
1p4
1o4
1i4
0K5
0I5
0D5
0C5
0B5
0=5
0<5
0;5
085
075
065
045
025
0I8
1F8
1D8
0B8
1>8
1=8
0:8
188
178
168
058
138
1/8
1-8
0+8
0m)
0k)
0i)
0h)
0g)
0f)
0b)
0a)
0`)
0_)
0[)
0Z)
0V)
0T)
0R)
0Q)
0P)
0O)
0N)
0M)
0L)
0K)
1J)
0U,
1S,
1R,
1P,
1N,
1L,
1K,
0J,
1G,
1F,
1D,
1?,
0=,
0<,
1;,
19,
17,
15,
14,
13,
02,
0-,
0,,
0*,
0(,
0',
0&,
0%,
0!,
0~+
0}+
0|+
0x+
0w+
0s+
0q+
0o+
0n+
0m+
0l+
0k+
1j+
1O2
1N2
1M2
1L2
1K2
1I2
1H2
1F2
1E2
1D2
1C2
1A2
1@2
1?2
1>2
1<2
1;2
182
172
162
152
142
122
112
102
1/2
0.2
1w2
0u2
0s2
0q2
0p2
0o2
0n2
0j2
0i2
0h2
0g2
0c2
0b2
0^2
0\2
0Z2
0Y2
0X2
0W2
0V2
0U2
1T2
0#8
0!8
0}7
0|7
0{7
0z7
0v7
0u7
0t7
0s7
0o7
0n7
0j7
0h7
0f7
0e7
0d7
0c7
0b7
0a7
1`7
0#:
1":
1!:
1}9
1v9
0u9
0t9
1r9
1o9
0m9
0l9
1j9
0i9
1h9
1f9
1d9
0c9
0b9
0K:
0G:
0E:
0D:
0>:
07:
15:
02:
11:
00:
0.:
0-:
0,:
1*:
057
0/7
1.7
0-7
1+7
0(7
0'7
0~6
0}6
1|6
1{6
0z6
0y6
0x6
0v6
1u6
0t6
144
0,4
0)4
0'4
0%4
0$4
1#4
0"4
1!4
1~3
1|3
1{3
0z3
0o3
1n3
1[4
1Z4
1T4
1Q4
1O4
1M4
1L4
0K4
1J4
0F4
1D4
1C4
0:4
061
141
131
021
1-1
0*1
1)1
1$1
1#1
1~0
0}0
0{0
0y0
0u0
0\1
1Z1
0W1
0U1
1S1
1R1
0Q1
0P1
0O1
1M1
0K1
0J1
1C1
0@1
1?1
08.
0/.
1..
0+.
0*.
0&.
1$.
1#.
0~-
0|-
1w-
0u-
1t-
0a.
1_.
1W.
0V.
0U.
1S.
1R.
0I.
1F.
0A.
1@.
1?.
0>.
0?+
0>+
0=+
0;+
0:+
07+
04+
03+
00+
0++
0)+
0(+
0'+
0&+
0$+
0#+
0"+
0!+
0~*
0}*
0|*
0e+
0`+
0Z+
0Y+
0S+
0R+
0N+
0I+
1B+
#99000
1"
1T!
b0 N:
b100000000000000000000000000000000000 O:
b110111000010101100011000110110000100000 P:
b1100111100010011100111001001111010000 Q:
b1001000110101011111000110001011101100001 R:
b110001010001000110001100100010010000 S:
b1001100101000111110100101001011010011000 T:
b11010111000001011010110100101110100 U:
b1010100001000001100100001000010010000000 V:
b1110101100111010001011100111100000 X:
b1110001010001000101010100010000010000 Y:
b101100011001111010100001101101110011110 "F
b10010011100110010101001110010010000100000 #F
b1011010101001001010110101101111000111101001 $F
b100100101000110010101001010010000101000000000 %F
b10000001100000111100110111010010111101000001 &F
b111110010101000010101000101100000000000000 'F
b101111000100001101110011100111011011000000011110100001 xK
b100000100100010000000101011011100000010000 yK
b1001111101011000010010011100001001010111011101000000000 zK
b100000000100101110100110011010110101000100000000000000 {K
b1111100111101101111111010111010101101010001010000100100011101100 HQ
b10000000101001001010001000110000100010000000000000 IQ
b1111101111101010110000010000000100100000110101101101000000000000 P!
b1111111001010110011100100100011101010001101101010000110011011110 Q!
b1111111010011000001010001110010110000000010110111011111000001 R!
b1111100111110010000000101001101001111011101011001000100011101100 S!
b11000000001110110010001010000000 H!
b10110001111011110110001001100011 J!
b10010110101010110101100000101101 L!
b101110010110000100100101011100 N!
b10000011001000010000100100000 I!
b101011100111000011100001010 K!
b10110010101001110010011001100101 M!
b11011110100011100010100010111101 O!
0iY
1hY
1gY
1fY
1eY
0aY
0`Y
1^Y
0]Y
0\Y
0[Y
0XY
1WY
0VY
1UY
1TY
1RY
1QY
0LY
1KY
0JY
1IY
1HY
0FY
0EY
1CY
0AY
1@Y
0?Y
1=Y
1<Y
1;Y
09Y
17Y
02Y
01Y
1,Y
1+Y
1*Y
1a
1^
1]
0Y
1X
0U
1T
0S
1Q
1P
0M
1K
1J
0I
1H
1E
0D
1B
1?
0=
1<
09
07
06
05
01
00
1.
1,
1(
1'
1&
1%
1$
0JN
1IN
0FN
1EN
1CN
1@N
1>N
0=N
1;N
0:N
18N
17N
05N
14N
12N
11N
0,N
0&N
1"N
1mM
1jM
1iM
1fM
1eM
0dM
0bM
1aM
0`M
0_M
0[M
1YM
0VM
0UM
1TM
0SM
0RM
0OM
1LM
1KM
1IM
0HM
1FM
1EM
1DM
0BM
0AM
1:M
04M
12M
1.M
0+M
0%M
0!M
1|L
0{L
0zL
1yL
0xL
0vL
0tL
1sL
1]L
0[L
0ZL
0WL
1UL
1TL
1SL
0QL
0PL
0ML
0LL
1KL
1JL
0FL
1DL
0AL
1@L
1>L
0=L
1;L
19L
08L
17L
05L
04L
03L
00L
0/L
1-L
1*L
1(L
0PJ
1MJ
1JJ
0IJ
0HJ
1FJ
0EJ
0AJ
0@J
0>J
1=J
19J
08J
13J
0#J
0"J
0!J
1}I
0|I
0wI
1vI
0uI
0rI
1qI
1pI
0nI
1mI
1lI
1hI
1gI
1fI
0eI
0dI
0cI
0bI
0aI
1`I
1_I
0^I
0YI
1LI
0KI
0II
0FI
0EI
1DI
0CI
1BI
0AI
0>I
1=I
0:I
04I
13I
02I
00I
1.I
1+I
1fG
0bG
1`G
0\G
1XG
1WG
1UG
1TG
1RG
0QG
1PG
1MG
0LG
1CG
0BG
1AG
1?G
0=G
0;G
09G
03G
11G
1,G
1)G
1&G
1$G
1!G
0|F
0yF
1xF
1wF
0uF
1tF
1sF
1oF
0nF
1lF
0^F
1]F
1\F
1[F
0YF
0TF
0QF
1PF
0NF
0LF
0KF
1FF
1EF
1DF
1CF
0BF
1?F
0>F
18F
05F
0$D
0~C
0|C
0{C
0uC
0nC
1lC
0iC
1hC
0gC
0eC
0dC
0cC
1aC
0UC
1TC
1SC
1QC
1JC
0IC
0HC
1FC
1CC
0AC
0@C
1>C
0=C
1<C
1:C
18C
07C
06C
0eB
0_B
1^B
0]B
1[B
0XB
0WB
0PB
0OB
1NB
1MB
0LB
0KB
0JB
0HB
1GB
0FB
1.@
1-@
1'@
1$@
1"@
1~?
1}?
0|?
1{?
0w?
1u?
1t?
0k?
1_?
0W?
0T?
0R?
0P?
0O?
1N?
0M?
1L?
1K?
1I?
1H?
0G?
0<?
1;?
03?
11?
0.?
0,?
1*?
1)?
0(?
0'?
0&?
1$?
0"?
0!?
1x>
0u>
1t>
0e>
1c>
1b>
0a>
1\>
0Y>
1X>
1S>
1R>
1O>
0N>
0L>
0J>
0F>
0D<
1B<
1:<
09<
08<
16<
15<
0,<
1)<
0$<
1#<
1"<
0!<
0w;
0n;
1m;
0j;
0i;
0e;
1c;
1b;
0_;
0];
1X;
0V;
1U;
0P;
0K;
0E;
0D;
0>;
0=;
09;
04;
1-;
0$;
0#;
0";
0~:
0}:
0z:
0w:
0v:
0s:
0n:
0l:
0k:
0j:
0i:
0g:
0f:
0e:
0d:
0c:
0b:
0a:
0MR
0LR
0KR
0JR
0GR
0DR
0BR
0@R
0=R
0;R
0:R
08R
05R
04R
03R
00R
0/R
0.R
0-R
0,R
0+R
1*R
0;=
04=
03=
0.=
0)=
1(=
1'=
0$=
0"=
0rR
0kR
1iR
0hR
1gR
0eR
1bR
0`R
1_R
0ZR
1YR
1UR
1TR
1QR
04>
12>
1*>
0)>
0(>
1&>
1%>
0z=
0r=
1p=
0o=
0sS
0qS
0oS
0nS
0kS
0jS
0iS
1eS
0dS
0cS
1`S
1_S
1^S
0]S
0\S
0ZS
0XS
0WS
1SS
10A
1)A
0%A
1$A
1#A
0~@
1}@
0|@
1{@
1x@
1w@
0u@
0>T
1<T
1;T
06T
05T
13T
02T
01T
00T
0/T
1*T
1(T
0&T
1%T
1$T
1xS
1'B
1~A
0wA
1uA
1tA
0kA
0EU
0?U
1>U
0=U
1;U
08U
07U
00U
0/U
1.U
1-U
0,U
0+U
0*U
0(U
1'U
0&U
1~D
1{D
1wD
1pD
0oD
1nD
1mD
1lD
1gD
0fD
1bD
1`D
1^D
0hU
0gU
0fU
1eU
1dU
1cU
0bU
0aU
0\U
1ZU
0XU
1UU
1TU
0SU
1PU
0MU
0LU
1KU
1HU
1GU
0pE
1`E
0]E
0YE
0XE
0WE
1UE
0GH
1FH
1EH
1DH
1CH
0BH
1AH
0?H
0=H
1<H
1;H
1:H
19H
17H
16H
10H
0/H
0.H
1,H
1+H
0(H
0~G
1zG
0yG
1xG
1vG
0tG
0rG
0pG
0zH
1vH
0rH
0qH
1pH
0nH
0lH
1hH
1fH
1eH
1dH
0bH
1`H
1_H
0^H
1]H
1XH
05K
04K
03K
01K
0-K
1,K
0+K
1*K
0(K
1$K
0#K
0!K
1~J
1{J
1zJ
0yJ
1wJ
1vJ
1uJ
0sJ
0qJ
0nJ
1jJ
1iJ
1lK
0iK
0eK
1dK
0cK
1bK
0aK
0`K
1_K
0^K
1]K
0[K
1ZK
0WK
1VK
0TK
0PK
0NK
1IK
0BK
1$W
0"W
0!W
0}V
0|V
1zV
1yV
1xV
0wV
1vV
1rV
1pV
0oV
0nV
0kV
1iV
1hV
0fV
0eV
1dV
1cV
0bV
1aV
1_V
1\V
1[V
0ZV
0UV
0TV
1RV
1OV
1MV
1GQ
1?Q
1>Q
1=Q
0;Q
07Q
15Q
11Q
1.Q
0*Q
1(Q
0'Q
1#Q
0"Q
1!Q
0|P
0{P
0yP
0xP
1uP
1rP
1pP
1RW
1OW
1NW
0MW
0LW
1KW
1JW
0HW
0GW
0EW
1DW
0CW
1AW
1=W
19W
15W
01W
10W
0/W
0.W
0-W
1+W
1*W
0'W
0&W
0%W
0lO
1kO
0hO
1gO
1eO
1`O
0_O
1]O
0\O
1YO
1VO
1TO
1dP
1\P
1[P
1ZP
0XP
0TP
1RP
1NP
1KP
0GP
1EP
0DP
1@P
0?P
1>P
0;P
0:P
08P
07P
14P
11P
1/P
1FX
0DX
0CX
0AX
0@X
1>X
1=X
1<X
0;X
1:X
16X
03X
12X
11X
00X
1.X
1(X
1~W
1|W
1yW
1wW
1vW
1uW
0tW
1pW
0nW
0mW
1kW
1jW
0gW
0fW
0eW
0GQ
1BQ
0?Q
0>Q
0=Q
14Q
03Q
0+Q
1*Q
0(Q
1&Q
0$Q
0}P
0wP
0uP
0pP
1QD
1ND
1JD
1CD
0BD
1AD
1@D
1?D
1:D
09D
15D
13D
11D
0?V
09V
18V
07V
06V
04V
13V
10V
0/V
0)V
1'V
0%V
0$V
1#V
1~U
1|U
0yU
1xU
1wU
1tU
1sU
0~D
0{D
0xD
0wD
0pD
0nD
0mD
0lD
0jD
0hD
0gD
1^@
1W@
0S@
1R@
1Q@
0N@
1M@
0L@
1K@
1H@
1G@
0E@
0sT
0qT
0oT
0nT
1mT
0iT
0cT
0bT
0aT
1]T
0\T
0ZT
1YT
1XT
0UT
1TT
1IT
14A
11A
1-A
0,A
0(A
0'A
0#A
0!A
1~@
0}@
0{@
0y@
0m<
0f<
0e<
0`<
0[<
1Z<
1Y<
0V<
0T<
0ES
0DS
0CS
0BS
1<S
0:S
16S
14S
13S
00S
1/S
0+S
1(S
1%S
1$S
0#S
1!S
1|R
0:=
05=
0-=
0(=
0'=
0#=
0|<
1{<
0l<
0g<
0_<
0Z<
0Y<
0U<
0P<
1O<
0k=
0j=
0i=
0h=
0e=
1b=
0`=
0^=
0]=
1\=
1Z=
1Y=
0X=
0V=
1U=
0S=
0R=
1L=
1K=
1J=
0I=
1G=
1D=
0/>
1->
0'>
0&>
0">
1}=
0w=
0v=
0u=
1t=
1b@
1_@
1[@
0Z@
0V@
0U@
0Q@
0O@
1N@
0M@
0K@
0I@
0eA
0cA
0aA
0`A
1_A
1^A
0[A
0WA
1UA
0TA
0RA
0QA
0OA
0MA
0JA
1HA
1FA
0EA
1;A
00B
1,B
1(B
0&B
1%B
1#B
1"B
1|A
1zA
1yA
0uA
0QD
0ND
0KD
0JD
0CD
0AD
0@D
0?D
0=D
0;D
0:D
0SE
0ME
1LE
0JE
1GE
0CE
0<E
1:E
08E
07E
13E
12E
1.E
1+E
1*E
1)E
1tE
1pE
1gE
1dE
1cE
0_E
0ZE
1YE
0VE
0UE
0dP
1_P
0\P
0[P
0ZP
1QP
0PP
0HP
1GP
0EP
1CP
0AP
0<P
06P
04P
0/P
1CO
1BO
0AO
0@O
0>O
0=O
1;O
17O
16O
13O
12O
1/O
0.O
1-O
1,O
1+O
1)O
0#O
1"O
0|N
1zN
0yN
0wN
0rN
0qN
1pN
0jN
1hN
1gN
0dN
0cN
0bN
1zO
1yO
0vO
0rO
1nO
0mO
0kO
0eO
1cO
0bO
1^O
0]O
1[O
0VO
1SO
1OO
1MO
1DO
0BO
1=O
1:O
19O
08O
0/O
1.O
0&O
0%O
1#O
0!O
0}N
1xN
1rN
0pN
0kN
0zO
0yO
1oO
0nO
1eO
0cO
1aO
0ZO
0TO
0KE
0HE
1EE
1DE
0=E
1;E
0:E
09E
17E
15E
14E
0qE
0pE
0gE
0cE
0aE
0`E
0bA
0_A
1[A
0ZA
0VA
0UA
1QA
1OA
1NA
1MA
1KA
1IA
13B
10B
0"B
0~A
0|A
0zA
0xA
0d=
1_=
1W=
1R=
0Q=
0M=
0H=
0G=
0,>
0$>
0}=
1r=
#100800
b1010101011110000100010110101010 d
b11001110110011001100110010011101 e
0"
1)Y
1'Y
1&Y
1%Y
0$Y
1"Y
0!Y
1}X
1|X
0zX
1yX
1xX
1tX
0rX
1pX
1nX
1mX
1lX
0kX
1iX
1hX
1u!
1s!
1r!
1q!
0p!
1n!
0m!
1k!
1j!
0h!
1g!
1f!
1b!
0`!
1^!
1\!
1[!
1Z!
0Y!
1W!
1V!
1fX
1dX
1bX
1_X
0^X
1]X
0ZX
1YX
0WX
0VX
1QX
1OX
1MX
1KX
0HX
1F!
1A!
1?!
1:!
09!
08!
14!
12!
01!
1/!
1+!
0*!
1(!
0'!
1%!
1$!
1~
0}
1|
1x
0r
1q
0p
0o
1k
0i
0T!
1r(
1p(
1o(
1n(
0m(
1k(
0j(
1h(
1g(
0e(
1d(
1c(
1_(
0](
1[(
1Y(
1X(
1W(
0V(
1T(
1S(
16"
14"
12"
1/"
0."
1-"
0*"
1)"
0'"
0&"
1!"
1}!
1{!
1y!
0v!
b0 yQ
b0 dQ
b0 ^Q
b0 XQ
b1 RQ
b1 LQ
b1 OQ
1VQ
0\Q
1_Q
0bQ
1eQ
1hQ
0nQ
0qQ
0tQ
0wQ
b1100010011001100110011011000101 KQ
b110001001100110011001101100010 NQ
b110001001100110011001101100010 QQ
b110001001100110011001101100010 TQ
b110011101100110011001100100111010 WQ
b111001110110011001100110010011101 ZQ
b0 ]Q
b111001110110011001100110010011101 `Q
b0 cQ
b1100010011001100110011011000101 fQ
b110011101100110011001100100111010 lQ
b111001110110011001100110010011101 oQ
b111001110110011001100110010011101 rQ
b111001110110011001100110010011101 uQ
b111001110110011001100110010011101 xQ
1")
0~(
1}(
0|(
1{(
1z(
0x(
0w(
0v(
0u(
0p'
0k'
0h'
0e'
0a'
0`'
1_'
0]'
1['
0Y'
0T'
1P'
1N'
1M'
1L'
1I'
1F'
1E'
1B'
1A'
1>'
1='
1:'
19'
17'
16'
15'
12'
11'
10'
1/'
1-'
1,'
1+'
1('
1%'
1$'
1!'
1~&
1{&
1z&
1w&
1v&
1t&
1s&
1r&
1o&
1n&
1m&
1l&
1j&
1i&
1h&
1e&
1b&
1a&
1^&
1]&
1Z&
1Y&
1V&
1U&
1S&
1R&
1Q&
1N&
1M&
1L&
1J&
1H&
1G&
1@&
1?&
0>&
1<&
1;&
09&
18&
17&
06&
05&
14&
13&
11&
10&
1,&
1+&
0f%
0d%
0c%
0\%
0[%
1Z%
0X%
0W%
1U%
0T%
0S%
1R%
1Q%
0P%
0O%
0M%
0L%
0H%
0G%
0F%
0E%
0D%
0C%
0B%
0@%
0?%
0=%
0<%
0;%
0:%
08%
07%
06%
05%
03%
02%
0/%
0.%
0-%
0,%
0+%
0)%
0(%
0'%
0&%
1%%
1#%
1"%
1!%
0~$
1|$
0{$
1y$
1x$
0v$
1u$
1t$
1p$
0n$
1l$
1j$
1i$
1h$
0g$
1e$
1d$
1c$
0b$
0a$
0`$
0_$
0^$
0]$
0[$
0Z$
0X$
0W$
0V$
0U$
0S$
0R$
0Q$
0P$
0N$
0M$
0J$
0I$
0H$
0G$
0F$
0D$
0C$
0B$
1A$
1?$
1>$
1=$
0<$
1:$
09$
17$
16$
04$
13$
12$
1.$
0,$
1*$
1($
1'$
1&$
0%$
1#$
1"$
1!$
0~#
0|#
1y#
0x#
0w#
1v#
0u#
0t#
0p#
0m#
0e#
1b#
0a#
0`#
0]#
0[#
0Z#
0Y#
1W#
0V#
1T#
0S#
0R#
0N#
0K#
0D#
0C#
0B#
1@#
0?#
0>#
0=#
1;#
17#
16#
14#
13#
10#
1/#
1,#
1+#
1(#
1'#
1$#
1~"
1}"
1x"
1t"
1s"
1q"
1p"
1m"
1l"
1i"
1h"
1e"
1d"
1a"
1]"
1\"
1X"
1V"
1R"
1Q"
1O"
1N"
1K"
1J"
1G"
1F"
1C"
1B"
1?"
1;"
1:"
16(
14(
18(
0<(
0@(
0D(
0R(
0m8
1m)
1k)
1g)
1f)
1d)
1c)
1`)
1_)
1\)
1[)
1X)
1W)
1T)
1P)
1O)
13*
10*
1,*
1+*
1)*
1(*
1%*
1$*
1!*
1~)
1{)
1z)
1w)
1s)
1r)
1/,
1,,
1(,
1',
1%,
1$,
1!,
1~+
1{+
1z+
1w+
1v+
1s+
1o+
1n+
0y,
0w,
1t,
0s,
0r,
1q,
0p,
0o,
0k,
0h,
0`,
1],
0\,
0[,
0F8
0A8
0>8
0;8
078
068
158
038
118
0/8
0*8
1#8
1!8
1~7
1}7
1z7
1w7
1v7
1s7
1r7
1o7
1n7
1k7
1j7
1h7
1g7
1f7
1c7
1b7
1a7
0`7
1s5
1q5
1p5
1o5
1l5
1i5
1h5
1e5
1d5
1a5
1`5
1]5
1\5
1Z5
1Y5
1X5
1U5
1T5
1S5
0R5
1M5
1K5
1J5
1I5
1F5
1C5
1B5
1?5
1>5
1;5
1:5
175
165
145
135
125
1/5
1.5
1-5
0,5
1&5
1$5
1#5
1z4
1y4
0x4
1v4
1u4
0s4
1r4
1q4
0p4
0o4
1n4
1m4
1k4
1j4
1f4
1e4
0d4
0Q2
0N2
0L2
0K2
0D2
0C2
1B2
0@2
0?2
1=2
0<2
0;2
1:2
192
082
072
052
042
002
0/2
1.2
0)2
0(2
0'2
0&2
0%2
0#2
0"2
0~1
0}1
0|1
0{1
0y1
0x1
0w1
0v1
0t1
0s1
0p1
0o1
0n1
0m1
0l1
0j1
0i1
0h1
0g1
1f1
0y/
1w/
1u/
1t/
1s/
0r/
1p/
0o/
1m/
1l/
0j/
1i/
1h/
1d/
0b/
1`/
1^/
1]/
1\/
0[/
1Y/
1X/
1W/
0V/
0Q/
0P/
0O/
0N/
0M/
0L/
0J/
0I/
0G/
0F/
0E/
0D/
0B/
0A/
0@/
0?/
0=/
0</
09/
08/
07/
06/
05/
03/
02/
01/
10/
0-/
1+/
1)/
1(/
1'/
0&/
1$/
0#/
1!/
1~.
0|.
1{.
1z.
1v.
0t.
1r.
1p.
1o.
1n.
0m.
1k.
1j.
1i.
0h.
1U,
0S,
0Q,
0P,
0O,
1M,
0L,
1J,
0I,
0H,
0D,
0A,
0:,
09,
08,
16,
05,
04,
03,
12,
091
171
151
031
001
0)1
0(1
0$1
0#1
0"1
0!1
0~0
0z0
0w0
1u0
1q0
0p0
0]1
1[1
0Z1
1X1
0V1
1T1
0S1
0R1
1Q1
1P1
0N1
1L1
1H1
1D1
0C1
1A1
1@1
0?1
0>1
1<1
044
034
114
004
0.4
1,4
0+4
1*4
1)4
0(4
1%4
0#4
1"4
0~3
0}3
1x3
0w3
0u3
1t3
1s3
0q3
1p3
0]4
0Z4
0Y4
0W4
0T4
0R4
0Q4
0O4
0M4
0L4
0J4
0D4
0C4
0B4
0@4
0>4
0=4
127
117
107
1/7
0.7
1,7
0+7
1*7
1%7
1"7
1x6
1v6
0u6
1s6
1m6
0l6
1W7
1V7
1U7
1S7
1P7
1O7
1L7
1K7
1H7
1G7
1D7
1C7
1A7
1@7
1?7
1>7
1<7
1;7
197
1;.
19.
18.
17.
13.
00.
1/.
0-.
1,.
1+.
0).
1'.
0!.
1|-
1z-
0x-
0t-
0_.
0].
0[.
1Y.
1X.
0W.
1U.
0T.
0S.
1Q.
0O.
1I.
0F.
0D.
1B.
0@.
0?.
1>.
1?+
1>+
1;+
19+
18+
16+
14+
12+
10+
1.+
1,+
1*+
1(+
1'+
1$+
1"+
1e+
1^+
1[+
1W+
1S+
1O+
1G+
1%:
0!:
1|9
1{9
0y9
1t9
0o9
1l9
0k9
0j9
0h9
0e9
1c9
1b9
1G:
0C:
1A:
17:
13:
12:
10:
1-:
0*:
#102600
1"
1T!
b10100110101010101010101101001100 N:
b100001000000010001000100010010000001 O:
b100110010110001100110011011010100111101 P:
b10001101000110011001100100111010000000 Q:
b101010010001000000000000001010100110100 R:
b10001100110011001100110010001001000000 S:
b1010111000100110011001100110110001000000 T:
b10000 U:
b110100100101001100110011000101001111000 V:
b1011011110110011001100110010111000000 W:
b111010000010101010101010111110100100 X:
b1010101111101010101010101000001010000 Y:
b10100011101000101101011010010111000000000 "F
b1010100000010010000100001001000010000000 #F
b1001011010011110101110100000001011010000000001 $F
b100101100001010101011101110010101001000000 %F
b11110011101111110001000111001111010010000000 &F
b100000000001010101000100000100000000000 'F
b101101010000101110001111100111011110111101011011110 xK
b100100101011000111010100001100100100000000 yK
b1111110100001111001110101010000010100110000001000000000 zK
b10100000110001010101101001010000000100000000000 {K
b1111100101100111110101100001100001111111010110111011111000001 HQ
b1000000001010011000001010010110011010000000100000000000000000000 IQ
b1110111110010010111000101000110010010001101111100011000101000010 P!
b1111101111101010110000010000000100100000110101101101000000000000 Q!
b1111111001010110011100100100011101010001101101010000110011011110 R!
b1111111010011000001010001110010110000000010110111011111000001 S!
b1010101011110000100010110101010 H!
b11000000001110110010001010000000 J!
b10110001111011110110001001100011 L!
b10010110101010110101100000101101 N!
b11001110110011001100110010011101 I!
b10000011001000010000100100000 K!
b101011100111000011100001010 M!
b10110010101001110010011001100101 O!
0hY
0gY
0fY
0eY
0cY
0bY
0_Y
0^Y
1]Y
1[Y
1ZY
0YY
1XY
0TY
1SY
0QY
0MY
1LY
0KY
0HY
0GY
0CY
1AY
0@Y
0=Y
0<Y
1:Y
07Y
16Y
05Y
14Y
12Y
11Y
0/Y
1c
0a
0`
0^
1[
1Z
1Y
0X
1W
1V
1U
0T
1S
1R
0Q
0N
0L
0K
0J
0H
0E
1D
0B
1A
0<
1;
0:
19
13
0.
1*
1)
0&
0%
0$
1LN
0IN
0EN
1DN
0CN
1BN
0AN
0@N
1?N
0>N
1=N
0;N
1:N
07N
16N
04N
00N
0.N
1)N
0"N
0kM
0jM
0iM
0gM
0cM
1bM
0aM
1`M
0^M
1ZM
0YM
0WM
1VM
1SM
1RM
0QM
1OM
1NM
1MM
0KM
0IM
0FM
1BM
1AM
0:M
16M
02M
01M
10M
0.M
0,M
1(M
1&M
1%M
1$M
0"M
1~L
1}L
0|L
1{L
1vL
0]L
1\L
1[L
1ZL
1YL
0XL
1WL
0UL
0SL
1RL
1QL
1PL
1OL
1ML
1LL
1FL
0EL
0DL
1BL
1AL
0>L
06L
12L
01L
10L
1.L
0,L
0*L
0(L
1PJ
0MJ
0LJ
1@J
0=J
0;J
09J
06J
04J
03J
02J
0%J
0}I
1|I
0{I
0zI
0xI
1wI
1uI
1tI
0sI
0mI
0lI
1kI
0iI
0hI
1eI
1dI
1cI
1bI
1^I
1[I
1ZI
1YI
1QI
1JI
1FI
1EI
0DI
1CI
1AI
19I
08I
07I
14I
0+I
0cG
0aG
0`G
0_G
0^G
1\G
0XG
0UG
0TG
0RG
0PG
1LG
1IG
0HG
1GG
1FG
1DG
0CG
19G
01G
1/G
0,G
1*G
0)G
1'G
0&G
0%G
0$G
1"G
0!G
0}F
0wF
0tF
0sF
0rF
1qF
1mF
0lF
0]F
0\F
0[F
0ZF
0WF
0VF
1TF
0RF
1QF
0PF
0OF
1NF
1LF
1KF
0JF
1IF
0HF
1GF
0EF
0CF
0?F
1>F
1=F
1<F
0;F
0:F
16F
1~C
0zC
1xC
1nC
1jC
1iC
1gC
1dC
0aC
1WC
0SC
1PC
1OC
0MC
1HC
0CC
1@C
0?C
0>C
0<C
09C
17C
16C
1,C
1+C
1*C
1(C
1%C
1$C
1!C
1~B
1{B
1zB
1wB
1vB
1tB
1sB
1rB
1qB
1oB
1nB
1lB
1bB
1aB
1`B
1_B
0^B
1\B
0[B
1ZB
1UB
1RB
1JB
1HB
0GB
1EB
1?B
0>B
00@
0-@
0,@
0*@
0'@
0%@
0$@
0"@
0~?
0}?
0{?
0u?
0t?
0s?
0q?
0o?
0n?
0_?
0^?
1\?
0[?
0Y?
1W?
0V?
1U?
1T?
0S?
1P?
0N?
1M?
0K?
0J?
1E?
0D?
0B?
1A?
1@?
0>?
1=?
04?
12?
01?
1/?
0-?
1+?
0*?
0)?
1(?
1'?
0%?
1#?
1}>
1y>
0x>
1v>
1u>
0t>
0s>
1q>
0h>
1f>
1d>
0b>
0_>
0X>
0W>
0S>
0R>
0Q>
0P>
0O>
0K>
0H>
1F>
1B>
0A>
0B<
0@<
0><
1<<
1;<
0:<
18<
07<
06<
14<
02<
1,<
0)<
0'<
1%<
0#<
0"<
1!<
1z;
1x;
1w;
1v;
1r;
0o;
1n;
0l;
1k;
1j;
0h;
1f;
0`;
1];
1[;
0Y;
0U;
1P;
1I;
1F;
1B;
1>;
1:;
12;
1$;
1#;
1~:
1|:
1{:
1y:
1w:
1u:
1s:
1q:
1o:
1m:
1k:
1j:
1g:
1e:
1MR
1LR
1KR
1HR
1ER
1AR
1=R
19R
15R
14R
11R
1?=
1>=
1;=
19=
18=
16=
14=
12=
10=
1.=
1,=
1*=
1(=
1'=
1$=
1"=
1wR
1uR
1tR
1sR
1rR
0pR
0oR
0nR
1jR
0iR
0fR
1eR
0dR
1cR
0bR
1]R
1\R
1ZR
0YR
0XR
0WR
1VR
0UR
0SR
0QR
02>
1+>
0*>
1(>
1z=
1s=
0p=
0vS
1tS
1rS
1qS
0pS
1oS
1nS
0mS
0lS
1jS
1hS
0gS
1dS
0bS
1aS
0_S
0^S
1]S
1\S
1YS
1XS
1WS
0VS
1US
0SS
1RS
0OS
17A
15A
00A
0/A
0*A
0)A
1(A
1%A
0$A
1!A
0~@
1|@
0z@
1u@
1t@
1q@
1p@
0=T
16T
14T
10T
1/T
0.T
1,T
1+T
0*T
0)T
0%T
1~S
1|S
0{S
1zS
0,B
0'B
0%B
0$B
0}A
0{A
0tA
0sA
0qA
0nA
1BU
1AU
1@U
1?U
1=U
0;U
17U
06U
15U
13U
1/U
0.U
1+U
1&U
1#U
0"U
0~T
1}T
0|T
1$E
1#E
1"E
1!E
1|D
1zD
1vD
1uD
1rD
1nD
1jD
1hD
1eD
0bD
1_D
1iU
0eU
0dU
1bU
1aU
1`U
0_U
0^U
0ZU
0UU
0TU
0RU
0QU
1OU
1NU
1MU
0KU
0JU
1IU
0HU
0GU
0nE
1]E
1[E
1XE
0FH
0EH
0DH
0CH
0AH
0@H
1=H
0;H
0:H
09H
07H
06H
05H
13H
01H
00H
1/H
0-H
0,H
0+H
1(H
1'H
0%H
1"H
0!H
1~G
1}G
1|G
1{G
0zG
1pG
0sH
1qH
0pH
0oH
1nH
1lH
0jH
1iH
0hH
1gH
0fH
0eH
0`H
0_H
1\H
0[H
1VH
0UH
1:K
15K
13K
1'K
0"K
1!K
0~J
1}J
0|J
1yJ
1xJ
0wJ
0uJ
1sJ
1rJ
1pJ
1nJ
0mJ
0lK
1eK
0dK
1`K
0\K
1YK
0XK
0VK
1TK
0RK
0QK
1PK
1NK
0KK
0IK
0$W
1#W
1"W
1!W
1~V
1|V
0zV
0yV
0xV
1wV
0vV
1sV
0rV
1oV
0jV
0hV
1fV
1eV
1bV
0aV
0`V
1WV
0VV
1UV
1SV
0QV
0OV
0MV
1FQ
1EQ
1DQ
1CQ
0BQ
1AQ
1<Q
01Q
10Q
0/Q
1,Q
1+Q
0)Q
1(Q
0&Q
0!Q
1zP
1yP
1xP
1vP
1uP
1tP
1sP
0PW
0NW
0DW
1BW
0AW
1@W
0?W
0=W
0<W
0;W
0:W
09W
18W
06W
04W
12W
11W
00W
1.W
0,W
0+W
1'W
1&W
1%W
0gO
1fO
0`O
1_O
1\O
0YO
0RO
0DO
1cP
1bP
1aP
1`P
0_P
1^P
1YP
0NP
1MP
0LP
1IP
1HP
0FP
1EP
0CP
0>P
19P
18P
17P
15P
14P
13P
12P
0FX
1EX
1DX
1CX
1BX
1@X
0>X
0=X
0<X
1;X
0:X
17X
06X
13X
02X
10X
0.X
1,X
1*X
1)X
0%X
1#X
1"X
0!X
1}W
0|W
0{W
1zW
0wW
0vW
0uW
1tW
1sW
0rW
0pW
0oW
1nW
0lW
0kW
1gW
1fW
1eW
0FQ
0EQ
0DQ
0CQ
0AQ
1>Q
0<Q
1;Q
17Q
04Q
0+Q
1%Q
0yP
0vP
0tP
0rP
1UD
1TD
1SD
1RD
1OD
1MD
1ID
1HD
1ED
1AD
1=D
1;D
18D
05D
12D
1<V
1;V
1:V
19V
05V
03V
02V
01V
1.V
0,V
1)V
1%V
0#V
0"V
0}U
1yU
0xU
1uU
0tU
0sU
0$E
0#E
0"E
0!E
1}D
1wD
1fD
1bD
0_D
0^D
1e@
1c@
0^@
0]@
0X@
0W@
1V@
1S@
0R@
1O@
0N@
1L@
0J@
1E@
1D@
1A@
1@@
0vT
1tT
1rT
1qT
0pT
1oT
1nT
0mT
0jT
1hT
0gT
0eT
1dT
1cT
1bT
1aT
1\T
0[T
1ZT
0WT
1VT
1UT
0TT
1ST
1RT
1MT
0LT
1KT
07A
05A
04A
01A
1/A
0%A
0"A
0!A
0w@
0t@
0s@
0p@
1q<
1p<
1m<
1k<
1j<
1h<
1f<
1d<
1b<
1`<
1^<
1\<
1Z<
1Y<
1V<
1T<
1ES
1CS
1BS
1AS
1?S
0<S
0;S
09S
17S
06S
15S
03S
12S
10S
0/S
1-S
0,S
1*S
1'S
0&S
0%S
0$S
1#S
1"S
0~R
0|R
0>=
08=
04=
0$=
0p<
0j<
0f<
0V<
1k=
1g=
0c=
0a=
1`=
0_=
1^=
1]=
1[=
0Z=
0Y=
0U=
0T=
1S=
1Q=
1P=
0N=
1M=
0K=
0J=
1I=
1H=
0F=
0D=
16>
15>
12>
10>
1/>
1,>
0(>
1'>
1#>
1!>
0~=
0{=
1y=
1v=
0t=
0s=
1o=
0e@
0c@
0b@
0_@
1]@
0S@
0P@
0O@
0G@
0D@
0C@
0@@
0hA
1fA
1eA
1dA
1bA
1aA
1`A
1_A
0^A
1]A
0\A
1ZA
0YA
1XA
1UA
1TA
1RA
0OA
0MA
1JA
0IA
0HA
0GA
0FA
0AA
0@A
1?A
0>A
1=A
14B
03B
00B
0.B
0)B
0(B
1'B
1$B
0#B
1~A
1{A
0yA
1wA
1vA
1tA
1sA
1pA
1oA
0UD
0TD
0SD
0RD
1PD
1JD
19D
15D
02D
01D
1PE
0LE
0FE
0EE
1CE
0@E
0?E
1=E
0;E
19E
06E
05E
03E
02E
0.E
1,E
0+E
0*E
0)E
1{E
1zE
1yE
1xE
1rE
1nE
1lE
1kE
1gE
1bE
1aE
1^E
0[E
1ZE
1WE
1VE
0cP
0bP
0aP
0`P
0^P
1[P
0YP
1XP
1TP
0QP
0HP
1BP
08P
05P
03P
01P
0CO
1BO
1>O
0<O
0;O
0:O
09O
18O
14O
03O
00O
1/O
0-O
0,O
0*O
0)O
1$O
0#O
0"O
1!O
1~N
1}N
1|N
1yN
0xN
1wN
0uN
0rN
0nN
1mN
0lN
1kN
0iN
0hN
1dN
1cN
1bN
1#P
1"P
1!P
1|O
1pO
0oO
1mO
1iO
1gO
0dO
1cO
0aO
0_O
0\O
0[O
1ZO
1WO
1TO
1RO
1PO
0OO
0MO
1KO
1AO
1@O
1?O
0>O
1<O
19O
07O
06O
02O
0/O
1&O
0~N
0tN
1qN
0oN
0mN
0#P
0"P
0!P
0|O
1vO
1rO
0fO
1`O
0SO
1OE
1NE
1ME
1LE
1JE
0DE
13E
0/E
0,E
1+E
0{E
0zE
0yE
0xE
1pE
1[E
0WE
0eA
1cA
0bA
0_A
0]A
1SA
1PA
1OA
1GA
1DA
0CA
1@A
04B
1.B
0$B
0!B
0~A
0vA
0sA
0oA
1h=
0b=
0^=
1N=
05>
0y=
